  
    Generic Library       2         4�         4�    �         :         :    �         p�         p�    �         k         k    �         ��         ��    �                ��  T��O FFSRCTRL.CKT4 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\FFSRCTRL.CKT FFSRCTRL.CKTR 3n W�    S 3n W�   Ctrl  W�   Q rl  W�    No Q  W�   ����������  �� �� �� �� ��
  ������ : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&      : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     ������ : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     	 : Generic Library                                �          ,�         ,�    �      �?N ��     �?N ��   �   	        ��&          ��   	     ��                         ��            ��        	      ��  	         Generic Library         !                         �         J                             Generic Library                                   �        Ctrl                          Generic Library         !                         �         K                             Generic Library         I        �         �    �        Q                              Generic Library         I        ��         ��    �   
     no Q                          A Generic Library       ,                         �         ��         ��    �      �?N V�     �?N V�   �           ��-       A Generic Library       *                         �         ��         ��    �       �?N V�     �?N V�   �           ��-        Generic Library       <        v/         v/    �   	      �         �    �         �         �    �         ��         ��    �       $     	  ��  
��O FFD.CKT/ C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\FFD.CKT FFD.CKTD �< ��E    Ctrl  ��E   Q rl  ��E    No Q  ��E   ��������  �� �� �� ��
  �� = Generic Library                                �         ��         ��    �       ��)     �� : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&      : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     ������ : Generic Library                                 �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     	 : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �   	        ��&          ��                 	                      ��            ��        	      ��     	    	 = Generic Library       4                         �   	   �?N �%     �?N �%   �      %  ��)     ����
 
                                 	                                                                  	     	        $ !             #             	   
        "         	                  "       
     % !   #  # &  &  ��* '   (            G     	  
    G 
     	    (            +          F          (            *           I           	 D          
 I            2              2            4   	         *            1          ,           +          +          F           D            /           )          H          H      
    + 
         ,            1            2            /             :            :              <           ! <         	 " )         # 1          $ <          	 % 9   	       	 & 1         ������          J     Ctrl     K     Q     no Q  ����                    L ��      �?N                                                          