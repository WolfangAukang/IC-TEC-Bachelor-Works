 
 
    Generic Library	                vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �   	      .I         .I    �   
      ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 <_<_    A1 <_<_   B0 <_<_   B1 <_<_   Ctrl0 <_   Z0 l0 <_    Z1 l0 <_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	               vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 <_<_    A1 <_<_   B0 <_<_   B1 <_<_   Ctrl0 <_   Z0 l0 <_    Z1 l0 <_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	       % 
 	      vw         vw    �   
      %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 <_<_    A1 <_<_   B0 <_<_   B1 <_<_   Ctrl0 <_   Z0 l0 <_    Z1 l0 <_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library               ,          ,    �         <*         <*    �         �)         �)    �         �)         �)    �          ��                            Generic Library                                  �         \�         \�    �        Ctrl                          Generic Library         -        �          �     �         �         �    �         b         b    �                      �        Z                              Generic Library                                   �         B�         B�    �         ��         ��    �         ��         ��    �       A                             Generic Library          
                        �         B�         B�    �         ��         ��    �         ��         ��    �       B                             Generic Library                                  �         B�         B�    �         ��         ��    �         ��         ��    �       C                           	  Generic Library                                  �         B�         B�    �         ��         ��    �         ��         ��    �       D                                                                                                                      	           
                                                                  	         	        	        	                                                                                        	   	    
      
       	   
                                     
              
                            %                   
              	                 %           % 
        	 
   	 #            
 %          -                   %           	 
    # 
          	 
    #                                                                                                                    
                        	     	                                                                                   Ctrl     Z     A     B     C   	  D 	                         ( ��       �An                                                         