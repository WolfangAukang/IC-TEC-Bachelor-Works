      Generic Library                                   �    	    Reset                         Generic Library                                  �         Set                         �� : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �   	        ��&      : Generic Library                                �          ,�         ,�    �      �?N ��     �?N ��   �           ��&       Generic Library         2        �R         �R    �        Q                              Generic Library         2        �Z         �Z    �   
     No Q                                                                                  
                       	   
  	                 	          
         '           '                                ' 	         2            "           	         
   
 2            "                        '            	                 	              	             
   ��          Set  ��    Reset      Q     No Q                  2 _ ��     �?N                                                          