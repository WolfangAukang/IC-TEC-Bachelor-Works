 
 	    Generic Library                                   �        R                             Generic Library                                  �         S                           �� : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&      : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&       Generic Library         2        2�         2�    �        Q                              Generic Library         2        ��         ��    �   
     No Q                           Generic Library          
                        �        Ctrl                         : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     	 : Generic Library                                �          ,�         ,�    �      �?N ��     �?N ��   �   	        ��&               	                                                       	          	              
                       	   
                        	          	          
         '           '                                ' 	         2            "           	    	        
 2            "                        '            	             	                               
   ��                    	                        	            
                  	                             S  ��    R      Q     No Q     Ctrl                      L ��       �?N                                                          