      Generic Library                                   �          C                             Generic Library                                  �        B                             Generic Library                                  �        A                             Generic Library         %                         �        Y                              Generic Library         %                         �   	     X                             = Generic Library                                 �      �?N Rw     �?N Rw   �        ��)      A Generic Library                                �         N         N    �      �?N �M     �?N �M   �   
        ��-       A Generic Library                                �         N         N    �      �?N �M     �?N �M   �           ��-       ] Generic Library                                �         �         �    �      �?N :�     �?N :�   �           ��M       	 = Generic Library                                �        N Rw       N Rw   �        ��)     
 M Generic Library                                �   	      ��         ��    �         ��         ��    �           ��;       A Generic Library                                �         N         N    �   	   �?N �M     �?N �M   �           ��-      
 
                                                    
                    	         
                    	    	  
                            	          	   
 
                                                                        %            $                                                              	 %           
         
                            	            	                                                                	        
     	       
          	     
              
                                                                                             C      B     A     Y     X                     $ 0 �^       �?N                                                          