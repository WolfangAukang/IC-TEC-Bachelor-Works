      Generic Library                                   �          A0                            Generic Library          	                        �        A1                            Generic Library                                  �        A2                            Generic Library                                  �        Hab                           Generic Library         1                         �        S0                             Generic Library         1                         �        S1                             Generic Library         1                         �        S2                             Generic Library         1                         �        S3                             Generic Library         1  
                       �        S4                           	  Generic Library         1                         �   	   	  S5                           
  Generic Library         1                         �   
   
  S6                             Generic Library         1                          �        S7                             Generic Library                �         �    �         �w         �w    �         �r         �r    �         �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �                    ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0  O�o    A1  O�o   Hab  O�o   C b  O�o    U b  O�o   D b  O�o   T b  O�o   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��    Generic Library                �         �    �         �w         �w    �   	      �r         �r    �   
      �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �         4           ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0   O�o    A1   O�o   Hab  O�o   C b  O�o    U b  O�o   D b  O�o   T b  O�o   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��   = Generic Library                                �      �?N ��     �?N ��   �   !   0  ��)      A Generic Library                                �         �0         �0    �   	   �?N z0     �?N z0   �   #   1   2  ��-       A Generic Library                                �         �0         �0    �      �?N z0     �?N z0   �       3     ��-                                                                                                            	         
               	         
                       ' '                              	  " 
    ! "  " $  $ #     %    %  &   ' &   '   (  ( )  )       *  * +  + 	  , 
  - ,   -   .  . /   /  ! 0   " 4 2 #  5 $  3 % 1 5 &  5 6 6                          	     
                   #    1            1 	           1            1            1          
 	 1   	        
 1   
         1 !                                            
    '            '           '           '                                        $ &    '          
  '           '           '                                    
                                     
             !   !            "       	    #            $          % 1         & 0         ' 0         ( /         ) /         * 0         + 0         , /         - /         . .         / . !         0         !   1        %   2         "  	 3        $   4        "  	 5      % # &              A0      A1     A2     Hab     S0     S1     S2     S3     S4  	 	  S5 	 
 
  S6 
    S7                                 	 	  
 
      0 ��     �An                                                         