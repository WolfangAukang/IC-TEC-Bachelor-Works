      Generic Library                $          $     �         ��         ��    �         ��         ��    �         ��         ��    �         �         �    �                 ��  d][Q
 LIBROS.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\LIBROS.CKT
 LIBROS.CKTC xg W�    B xg W�   A xg W�   Y xg W�    X xg W�   ����������  �� �� �� �� ��  ���������� = Generic Library                                 �      �?N Rw     �?N Rw   �        ��)      A Generic Library                                �         N         N    �      �?N �M     �?N �M   �   
        ��-       A Generic Library                                �         N         N    �      �?N �M     �?N �M   �           ��-       ] Generic Library                                �         �         �    �      �?N :�     �?N :�   �           ��M       	 = Generic Library                                �        N Rw       N Rw   �        ��)     
 M Generic Library                                �   	      ��         ��    �         ��         ��    �           ��;       A Generic Library                                �         N         N    �   	   �?N �M     �?N �M   �           ��-      
 
    ��         ��            ��                     
          ��         	         
          ��        	    	  
         Generic Library                  ,X         ,X    �         T         T    �                      �    	     LIbros                       ` Generic Library               �B         �B    �         B�         B�    �         ��         ��    �          ��         ��    �         R�         R�    �         �         �    �             ��	                                    ` Generic Library               ��         ��    �         �         �    �         ��         ��    �         b�         b�    �           ��                            Generic Library                                  �         b�         b�    �        Palabras                                                                                                                                                                                                  ��                 ����          LIbros     Palabras            	 1 ��       �?N                                                          