 # "    Generic Library                                   �         A                             Generic Library                                  �   2     B                             Generic Library                                  �   J     C                            A Generic Library                                �         L         L    �         �N         �N    �   1         ��-       = Generic Library                                �         S         S    �   I     ��)      M Generic Library                                  �         �W         �W    �         rY         rY    �            ��;        Generic Library         %        2l         2l    �        Q                             D Generic Library        
                        �         �]         �]    �         �b         �b    �   	      ng         ng    �              ��0       = Generic Library        
                         �         ~z         ~z    �        ��)     	 = Generic Library                                �         B         B    �   0     ��)     
 = Generic Library                                �         ʈ         ʈ    �   K     ��)       Generic Library            	      &�         &�    �        R                              Generic Library                 ��         ��    �   /     S                              Generic Library                 ^�         ^�    �        T                             = Generic Library                                 �   
      >�         >�    �      >  ��)     �� A Generic Library        1                        �         .         .    �         �         �    �         E  ��-       M Generic Library        /                         �         *>         *>    �         n�         n�    �   F        ��;        Generic Library         " 0       
         
    �      	  Z                             = Generic Library        1                        �         �         �    �        ��)       Generic Library          #       j�         j�    �   ,   
  X                              Generic Library                 ��         ��    �   #     W                             D Generic Library        '                        �         <         <    �         �8         �8    �         �         �    �              ��0       = Generic Library                                �         �         �    �   G   $  ��)      A Generic Library                                �         2�         2�    �         ^�         ^�    �   &   $   #  ��-       = Generic Library                                 �         �I         �I    �   +   &  ��)      M Generic Library                                �          nn         nn    �         �         �    �   8   9   6  ��;        Generic Library                 f         f    �   6     U                             = Generic Library                                 �         JJ         JJ    �   :   8  ��)      = Generic Library                                �         "�         "�    �   =   ;  ��)      A Generic Library         
                       �         �$         �$    �         Hv         Hv    �   >   ;     ��-       = Generic Library        (                        �         �         �    �   %     ��)       = Generic Library        )                        �         �|         �|    �   !     ��)     ! = Generic Library        '                         �         P�         P�    �   4     ��)     "  Generic Library         # (                        �        Y                                	                         !             	     	                                         
                                                        	         
    	          
                                             !                             "                                                                        . .      C   ) C  H    	     F  * H   E  	  	  	 
 ) !     3 %  . D  A )  @ I  J @  * 4  5 *     B L  B 3  5 +  A K  7 9  " /  < 7  < :   <  ' 0   H  ? =   ( 1 ! 2 ( " ( ' # L G $ 7 5 % " ? & , B ' ' " (   ) - C * ? L + @ A , 3 D - D  M G                                           	     %                " 1              ����  �          2         	       	     ������ # )      "                                                           	               
                        	   *                      (    ��               4      -     )               2                (  !                                   (                    2             /         !  *        
   "       ' %   #                $                %  )          &                '      "  '   (      " !     )  *     
    *  (          +             ,  $       &   -  �    )   .  �       /            0    	        1             2         !   3  )      ,   4  (  !         5       $     6                7        $    8                9            :             ;               <            =            >               
 ?       % *   @        +   A       +    B  $    &     C  2     )    D  4    ,  -   E  3          F  0           G          #   H  /          I            J            K    
        L       *  #       ' 
 ;  | Pedro Henrique rodriguez de Oliveira 2013086585 Fundamentos de organizaci�n de computadoras Grupo 1 Operaciones aritmeticas        A      B     C     Q     R     S     T  �� "  Y " 	   Z  
   X     U     W                                 	 
  
 	      / R�       �An                                                         