 
 	    Generic Library                                   �        D                            = Generic Library                                �         ��         ��    �       ��)     �� : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&      : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �           ��&       Generic Library         2        |�         |�    �        Q                              Generic Library         2        Ҧ         Ҧ    �   
     No Q                           Generic Library          
                        �        Ctrl                         : Generic Library                                 �         ,�         ,�    �      �?N ��     �?N ��   �           ��&     	 : Generic Library                                �         ,�         ,�    �      �?N ��     �?N ��   �   	        ��&                             	                                             	             	            
                      	   
                 ��  	                      !     	          
         '           '                                ' 	         2                        	    	        
 2            "                        '            	             	       ��        
    ��                    	                        	            
                   	                                                                              ��      ����    D      Q     No Q     Ctrl                 L ��       �?N                                                          