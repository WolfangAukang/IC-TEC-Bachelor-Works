     ` Generic Library      	         �\         �\    �                      �         2         2    �         ��         ��    �          b�         b�    �         ��         ��    �         J�         J�    �         vo         vo    �       R  U      ��
                                              Generic Library                �         �    �         �         �    �         r�         r�    �         �8         �8    �         |A         |A    �         4         4    �         ,=         ,=    �         ޟ         ޟ    �         4E         4E    �   	       P          P    �   
      �O         �O    �         
)         
)    �            .         
  	    >  ;  ��  ��O
 DEC3X8.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC3X8.CKT
 DEC3X8.CKTA0 ;_�;_    A1 ;_�;_   A2 ;_�;_   Hab _�;_   S0  _�;_    S1  _�;_   S2  _�;_   S3  _�;_   S4  _�;_   S5  _�;_   S6  _�;_   S7  _�;_  	 ������������������������  �� �� �� �� �� �� �� ��
 �� �� �� ��  ������������������������  Generic Library                �         �    �         �w         �w    �         �r         �r    �         �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �                    ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0 i W�    A1 i W�   Hab  W�   C b  W�    U b  W�   D b  W�   T b  W�   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��    Generic Library                �         �    �         �w         �w    �   	      �r         �r    �   
      �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �         4           ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0   W�    A1   W�   Hab  W�   C b  W�    U b  W�   D b  W�   T b  W�   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��   = Generic Library                                �      �?N ��     �?N ��   �   !   0  ��)      A Generic Library                                �         �0         �0    �   	   �?N z0     �?N z0   �   #   1   2  ��-       A Generic Library                                �         �0         �0    �      �?N z0     �?N z0   �       3     ��-           ��             ��          ��            ��                       ��        ��       ��       ��  	         
      ��       ��       ��       ��              Generic Library                                  �   P     Hab                           Generic Library                  �         �    �         X�         X�    �         �#         �#    �         j#         j#    �         A                             Generic Library                �         �    �         �         �    �         r�         r�    �         �8         �8    �         |A         |A    �         4         4    �         ,=         ,=    �         ޟ         ޟ    �         4E         4E    �          P          P    �         �O         �O    �         
)         
)    �   f   `      I               F  H  ��  ��O
 DEC3X8.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC3X8.CKT
 DEC3X8.CKTA0  ���    A1  ���   A2  ���   Hab  ���   S0   ���    S1   ���   S2   ���   S3   ���   S4   ���   S5   ���   S6   ���   S7   ���  	 ������������������������  �� �� �� �� �� �� �� ��
 �� �� �� ��  ������������������������  Generic Library                �         �    �         �w         �w    �         �r         �r    �         �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �                    ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0 i W�    A1 i W�   Hab  W�   C b  W�    U b  W�   D b  W�   T b  W�   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��    Generic Library                �         �    �         �w         �w    �   	      �r         �r    �   
      �7         �7    �         V�         V�    �         ��         ��    �         :�         :�    �         4           ��  R�O
 DEC2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\DEC2X4.CKT
 DEC2X4.CKTA0   W�    A1   W�   Hab  W�   C b  W�    U b  W�   D b  W�   T b  W�   ��������������  �� �� ��	 ��
 �� �� �� 
 ������������ = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-      ��     ��   	              ��     
                 	             
               	          
                       ��           	      ��   
      ��        ��        ��   = Generic Library                                �      �?N ��     �?N ��   �   !   0  ��)      A Generic Library                                �         �0         �0    �   	   �?N z0     �?N z0   �   #   1   2  ��-       A Generic Library                                �         �0         �0    �      �?N z0     �?N z0   �       3     ��-           ��             ��          ��            ��                       ��        ��       ��       ��  	         
      ��       ��       ��       ��              Generic Library                                  �        Out0                           Generic Library          	                        �         Out1                           Generic Library                                  �   !     Out2                           Generic Library                                  �   "     Out3                         	  Generic Library                                  �   #     Out4                         
  Generic Library           	                       �   $     Out5                           Generic Library           
                       �   ?     Out6                           Generic Library                                  �   :   	  Out7                           Generic Library                                  �   '   
  Out8                           Generic Library          !                        �   (     Out9                           Generic Library          $                        �   )     Out10                          Generic Library          '                        �   *     Out11                          Generic Library          *                        �   +     Out12                          Generic Library          -                        �   ,     Out13                          Generic Library          0                        �   -     Out14                          Generic Library          3                        �   G     Out15                         A Generic Library                                �         z�         z�    �      �?N *�     �?N *�   �   Q        ��-       A Generic Library                                �         z�         z�    �      �?N *�     �?N *�   �      N   O  ��-       ` Generic Library      
         "o         "o    �         ^>         ^>    �         >         >    �         �=         �=    �          n=         n=    �         =         =    �         �<         �<    �         ~<         ~<    �   b  c  d  e  a   ��
                                             = Generic Library      
 	                        �      �?N ��     �?N ��   �   S  K  ��)                                                                                               	    	     
    
                                                                                                                                       H H       
 2  / !   1  0    1 /   0     2 3 	 3 " 
 4 #  5 4  	 5  6 $  7 6   7   I  = (  8 ?  F E  ;   > 9  & :  8 9   &   D  < %  % )   *  @    A   @   A B ! B + " C , # E  $  < % C D &  = '  - ( .  )  ' * H J + G J , O  - M N . S T / M P 0 L  1   2 M  3 K Q 4 V S 5 U T 6 R  7 V W 8 W X 9 X L :  Y ; Y  < Z  = \ ] >  [ ? Z [ @  \ A ]  B  ^ C ^ _ D b f E _ a F c ` G d  g e   	                         1         6 :   ��          @      !      G               (                  	 	           
  
           	                                         0     	      ;           <            A               B        	     2 1            >   ��  "     ,            )            &     !      $     "           #           $           1    # '            (                  
          !            "         	   #    	     
   $    
       	 %  %        &          '         )   (  "          )  %          *  (          +  +       !   ,  .       "   -  1       '   .  
      (   /          0          1  	        2  
        3       	   4      
    5          6         	 7         	 8         
 9         
 :            ;           <  !     $   =        &   >          
 ?           
 @  "        A  #         B  +      !   C  .    " %   D  $    %    E  %    #    F  %         G  4       +   H  &      *   I  "         J  4    + *   K         3   L 
     0 9   M 	     - / 2   N        -   O         ,   P 	        /   Q         3   R         6   S  	       4 .   T  	    5 .   U         5   V 	 	    4 7   W 	     7 8   X 
     8 9   Y  	    : ;   Z      < ?   [      > ?   \      @ =    ]      = A    ^      B C       _ 
     C E       `         F   a 
        E       b         D    c         F   d  !      G   e  "         f         D              A     Hab     Out0     Out1     Out2     Out3   	  Out4 	  
  Out5 
    Out6  	   Out7  
   Out8     Out9     Out10     Out11     Out12     Out13     Out14     Out15                                 	 	  
 
                        L ��      �An                                                         