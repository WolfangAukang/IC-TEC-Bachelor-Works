 
 
    Generic Library                                   �          A                             Generic Library                                  �        B                             Generic Library                                  �        C                             Generic Library                                  �        D                             Generic Library                                  �    	    Ctrl0                         Generic Library         (        t         t    �        Z                              Generic Library                                  �    	    Ctrl1                         Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA � $    B � $   Ctrl  $   Z rl  $    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  $    B rl  $   Ctrl  $   Z rl  $    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   	  Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �         
     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  $    B rl  $   Ctrl  $   Z rl  $    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   	 	                                                           	         	          	     	                     
                  	   
                          	                                                                            	          	  	                	            
   	           
  
  	                                                               	                   %   	          (                                                       	          
                                                                  A      B     C     D     Ctrl0     Z     Ctrl1                            L ��       �An                                                         