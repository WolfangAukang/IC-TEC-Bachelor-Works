   ��  Generic Library                                   �         A                             Generic Library                                  �         B                             Generic Library                                  �        C                             Generic Library                                  �   #     D                             Generic Library          
                        �        E                             Generic Library         .        �         �    �        L-Z                            Generic Library         '        F�         F�    �        L-Y                            Generic Library                  �         �    �        L-X                          	  Generic Library                 ֕         ֕    �        L-V                          
  Generic Library                 �         �    �   $   	  L-R                            Generic Library                  �         �    �   &   
  L-S                            Generic Library         '  
      f�         f�    �   *     L-T                            Generic Library         .  	      �         �    �   .     L-U                            Generic Library         .        ��         ��    �        L-Q                            Generic Library                             �         �         �    �         8�         8�    �         ��         ��    �         ��         ��    �         Ȧ         Ȧ    �         ��         ��    �         T         T    �         �         �    �   	      ��         ��    �   
      Ч         Ч    �         Db         Db    �         �G         �G    �         �I         �I    �         $�         $�    �         ��         ��    �         �H         �H    �         `�         `�    �         t         t    �         <�         <�    �         tZ         tZ    �         �;         �;    �         N;         N;    �         ��         ��    �         �         �    �                   >  9  8    6  5  4  $  1  -  )  (  %          
  	    ��  �lQ
 086585.CKTJ C:\USERS\LEEECHER\DROPBOX\TEC\CLASES\FUNDA(~1\CIRCUI~2\CIRCUI~1\086585.CKT
 086585.CKTA  UE�    B  UE�   C  UE�   D  UE�   E  UE�   L-Z  UE�    L-Y  UE�   L-X  UE�   L-V  UE�   L-U  UE�   L-T  UE�   L-S  UE�   L-R  UE�   L-Q  UE�   L-P  UE�	   L-O  UE�
   L-N  UE�  
 L-L  UE�   L-K  UE�   L-J  UE�   L-I  UE�   L-H  UE�   L-G  UE�   L-M  UE�  	 L-F  UE�   ��������������������������������������������������  �� �� �� �� �� �� �� �� ��+ ��8 ��; ��> ��H ��P ��` ��g ��| �� ��� ��� ��� ��� ��o ��� ��� ��������������������������������������������������������������������������������������������������������������������������������������������F M Generic Library       +                        �         �#         �#    �      �?N �     �?N �   �     �   �  ��;      G A Generic Library                               �         �[         �[    �   	   �?N Dj     �?N Dj   �   �   �   �  ��-      H A Generic Library        
                         �         X         X    �      �?N ��     �?N ��   �   �   �   �  ��-      I = Generic Library                               �      �?N ��     �?N ��   �   �   �  ��)     J = Generic Library                                 �   
   �?N J�     �?N J�   �     �  ��)     K = Generic Library        
                       �      �?N >     �?N >   �      ��)     L A Generic Library        
                       �         ��         ��    �      �?N >     �?N >   �        ��-      M M Generic Library       !                        �   	      ��         ��    �      �?N �C     �?N �C   �     �   �  ��;      N = Generic Library                               �      �?N B/     �?N B/   �   ^  	 ��)     O A Generic Library       & 
                       �         �o         �o    �      �?N �     �?N �   �     �    ��-      P A Generic Library                               �         �         �    �      �?N ��     �?N ��   �        ��-      Q ] Generic Library                               �         &1         &1    �      �?N �\     �?N �\   �        ��M       ����T M Generic Library       ! �                        �         N�         N�    �      �?N �f     �?N �f   �         ��;      U M Generic Library        �                        �         V.         V.    �      �?N ޜ     �?N ޜ   �   #  !  " ��;      V A Generic Library        �                        �         �         �    �      �?N p.     �?N p.   �   $  4   ��-      W = Generic Library                                �      �?N &U     �?N &U   �   &  ' ��)     X = Generic Library        �                        �      �?N *     �?N *   �   -  ( ��)     Y A Generic Library        �                        �          �          �    �      �?N n�     �?N n�   �   +    ) ��-      Z A Generic Library        �                        �         �%         �%    �      �?N f!     �?N f!   �   (  '  + ��-      [ = Generic Library        �                        �      �?N v�     �?N v�   �     0 ��)     \ ] Generic Library        �                        �         ��         ��    �      �?N ��     �?N ��   �   3  2  $ ��M       ] A Generic Library        �                        �         ��         ��    �      �?N >�     �?N >�   �   <  8   ��-      ����������c M Generic Library       ! �                        �         �r         �r    �      �?N �W     �?N �W   �   H  \  9 ��;      d M Generic Library        �                        �         ��         ��    �      �?N ��     �?N ��   �   I  Y  G ��;      e A Generic Library        �                        �         �1         �1    �       �?N N�     �?N N�   �   L  K  O ��-      f A Generic Library        �                         �   !      �W         �W    �      �?N F�     �?N F�   �   T  S  R ��-      g = Generic Library        �                        �   !   �?N ʎ     �?N ʎ   �   J  S ��)     h = Generic Library        �                        �   "   �?N ʎ     �?N ʎ   �   M  V ��)     i A Generic Library        � #                       �   "      �W         �W    �      �?N F�     �?N F�   �   ]  V  F ��-      j M Generic Library        � $                       �   %      �%         �%    �      �?N Z%     �?N Z%   �   ^  g  B ��;      k = Generic Library        � &                       �   %   �?N n�     �?N n�   �   a  ` ��)     l M Generic Library        �                        �         �         �    �   &   �?N ��     �?N ��   �   b  _  a ��;      m A Generic Library        �                        �         �1         �1    �   #   �?N N�     �?N N�   �     N  X ��-      n A Generic Library        � '                       �   (      �}         �}    �   $   �?N �1     �?N �1   �   l  h  [ ��-      ��p M Generic Library       ! � )                       �   *      R�         R�    �   +   �?N ��     �?N ��   �   t    p ��;      q A Generic Library        � ,                       �   -      �b         �b    �   *   �?N �
     �?N �
   �   u  y  s ��-      r ] Generic Library        �                        �         r�         r�    �   ,   �?N Z     �?N Z   �   x  w  r ��M       s = Generic Library        �                        �   -   �?N 2�     �?N 2�   �   
  | ��)     t M Generic Library        � .                       �   /      ��         ��    �   )   �?N 2^     �?N 2^   �   }  ~  o ��;      u A Generic Library        � 0                       �         2[         2[    �   /   �?N v     �?N v   �   �  �  � ��-      v A Generic Library        �                        �         F-         F-    �   0   �?N ��     �?N ��   �   �  �  � ��-      w = Generic Library        �                        �   1   �?N F     �?N F   �   �  � ��)     x A Generic Library        �                        �   1      2^         2^    �   .   �?N r     �?N r   �   �   �  � ��-      ��z = Generic Library        �                        �   2   �?N �     �?N �   �   �  � ��)     { ] Generic Library        �                        �         �         �    �   3   �?N fq     �?N fq   �   �  �  � ��M       | A Generic Library        � 2                       �   3      RX         RX    �   4   �?N �\     �?N �\   �   �  �  � ��-      } A Generic Library        �                        �         "�         "�    �   5   �?N �~     �?N �~   �   �  �  � ��-      ~ A Generic Library        �                        �   5      ��         ��    �   6   �?N &�     �?N &�   �   �  �  � ��-       M Generic Library        � 4                       �   6      n�         n�    �   7   �?N v�     �?N v�   �   �  �  � ��;      � A Generic Library       ! �                        �   7      (         (    �   8   �?N �;     �?N �;   �   �   �  � ��-      ��� A Generic Library        � 9                       �   :      �         �    �   ;   �?N ��     �?N ��   �   �  �  � ��-      � A Generic Library        �                        �         �         �    �   :   �?N 
�     �?N 
�   �     �  � ��-      � A Generic Library        �                        �         Z�         Z�    �   9   �?N jw     �?N jw   �   �  �  � ��-      � M Generic Library        � <                       �   =      �P         �P    �   >   �?N V�     �?N V�   �   �  �  � ��;      � G Generic Library       > � ?                       �   @      vD         vD    �   A      n         n    �   B      �T         �T    �   C      �H         �H    �   �  �  �  �  � ��3     ��� = Generic Library        �                        �   D   �?N ��     �?N ��   �   �  � ��)     � M Generic Library        �                        �         *�         *�    �   =   �?N ��     �?N ��   �     �  � ��;      � M Generic Library        � D                       �         b�         b�    �   <   �?N *,     �?N *,   �   �  �  � ��;      ��� = Generic Library        �                        �   E   �?N �S     �?N �S   �   �  � ��)     � M Generic Library       ! � F                       �   G      &@         &@    �   H   �?N ��     �?N ��   �   �  �  � ��;      � A Generic Library        �                        �   E      �y         �y    �   G   �?N Fk     �?N Fk   �      �  � ��-      � M Generic Library        � I                       �   J      ��         ��    �   F   �?N j�     �?N j�   �   �  �  � ��;      � A Generic Library        � K                       �         ��         ��    �   J   �?N 2�     �?N 2�   �   �  �  � ��-      � A Generic Library        �                        �         >�         >�    �   K   �?N ��     �?N ��   �   �  �  � ��-      � A Generic Library        � L                       �   M      �s         �s    �   I   �?N R�     �?N R�   �   �  �  � ��-      � = Generic Library        �                        �   M   �?N '     �?N '   �   �   � ��)     � ] Generic Library        �                        �         ^+         ^+    �   L   �?N �3     �?N �3   �   �  �  � ��M       � M Generic Library       & � N                       �   O      ��         ��    �   P   �?N �;     �?N �;   �   �  �  � ��;      � M Generic Library       ! � Q                       �   R                   �   O   �?N ��     �?N ��   �   �  �  � ��;      � M Generic Library       ! � S                       �   T      f\         f\    �   N   �?N 6k     �?N 6k   �   �  �  � ��;      ��� = Generic Library        �                        �   U   �?N >�     �?N >�   �   �   � ��)     � = Generic Library        �                        �   V   �?N J�     �?N J�   �   �  � ��)     � A Generic Library        � W                       �         &�         &�    �   Q   �?N ��     �?N ��   �   �  �   � ��-      � A Generic Library        �                        �         ��         ��    �   W   �?N �     �?N �   �   �  �  � ��-      � A Generic Library        � V                       �   U      ��         ��    �   X   �?N �     �?N �   �   �  �  � ��-      � ] Generic Library        �                        �         �         �    �   Y   �?N �:     �?N �:   �        ��M       � A Generic Library        � X                       �         &�         &�    �   R   �?N ��     �?N ��   �   �  �  � ��-      � = Generic Library        �                        �   Z   �?N �7     �?N �7   �     	 ��)     � A Generic Library        � Y                       �   Z      V�         V�    �   T   �?N V�     �?N V�   �        ��-      � A Generic Library        � [                       �   \      V�         V�    �   S   �?N V�     �?N V�   �        � ��-      � = Generic Library        �                        �   \   �?N �7     �?N �7   �      ��)     � = Generic Library        � ]                       �   [   �?N "N     �?N "N   �       ��)     � ] Generic Library        �                        �         �         �    �   ]   �?N �:     �?N �:   �   !  �    ��M       ��� M Generic Library       & � ^                       �   _      B         B    �   `   �?N �=     �?N �=   �   -     ��;      � M Generic Library       ! | a                       �   b      �w         �w    �   ^   �?N ��     �?N ��   �      "   ��;      ��� = Generic Library        u                        �   c   �?N (�     �?N (�   �   '  * ��)     � = Generic Library        s                        �   d   �?N �     �?N �   �   �   + ��)     � M Generic Library        q e                       �   f      Z�         Z�    �   g   �?N ��     �?N ��   �   /  4  & ��;      � M Generic Library        s d                       �   c      jF         jF    �   f   �?N Nl     �?N Nl   �   +  *  0 ��;      � = Generic Library        o                        �   h   �?N �f     �?N �f   �   1  2 ��)     � M Generic Library        o h                       �         >�         >�    �   e   �?N ��     �?N ��   �   2  )  , ��;      � = Generic Library        �                        �   i   �?N J�     �?N J�   �   �   8 ��)     � = Generic Library        �                        �   j   �?N �     �?N �   �   <  9 ��)     � A Generic Library        � j                       �   i      ��         ��    �   k   �?N �     �?N �   �   9  8  ; ��-      � A Generic Library        � k                       �         &�         &�    �   _   �?N ��     �?N ��   �   ;  ?   ��-      � A Generic Library         l                       �         &�         &�    �   b   �?N ��     �?N ��   �   E  �    ��-      � A Generic Library        ~                        �         ��         ��    �   l   �?N �     �?N �   �   F  B  E ��-      � M Generic Library       & a m                       �   n      ��         ��    �   o   �?N ��     �?N ��   �   c  Y  H ��;      � A Generic Library        y p                       �   q      Z_         Z_    �   a   �?N N�     �?N N�   �   I  K  J ��-      � = Generic Library        { r                       �   q   �?N ��     �?N ��   �   O  K ��)     � ] Generic Library        z                        �         ��         ��    �   r   �?N N�     �?N N�   �   �   P  O ��M       � = Generic Library        x                        �   p   �?N �      �?N �    �   R  U ��)     � = Generic Library        d                        �   s   �?N <&     �?N <&   �   �  Z ��)     � A Generic Library       ! e s                       �   t      ��         ��    �   n   �?N �$     �?N �$   �   X  [  \ ��-      � = Generic Library        ` u                       �   v   �?N vx     �?N vx   �   b  M ��)     � A Generic Library        ` v                       �         z�         z�    �   m   �?N �     �?N �   �   M  `  V ��-      � ] Generic Library        _                        �         ��         ��    �   u   �?N ڄ     �?N ڄ   �   f  �   b ��M       � ] Generic Library        f                        �         Z�         Z�    �   w   �?N >�     �?N >�   �   �  �   a ��M       � A Generic Library        W                        �   x      ��         ��    �   y   �?N ��     �?N ��   �   n  q  p ��-      � = Generic Library        Y                        �   x   �?N "9     �?N "9   �   v  q ��)     � M Generic Library        h w                       �   z      �4         �4    �   t   �?N ��     �?N ��   �   +  �  r ��;      � A Generic Library        [                        �         n�         n�    �   {   �?N �     �?N �   �   �   x  w ��-      � A Generic Library        Y y                       �   {      �V         �V    �   |   �?N �R     �?N �R   �   |  {  z ��-      ����� A Generic Library        P }                       �   ~      �V         �V    �      �?N �R     �?N �R   �   �  �  ~ ��-      � A Generic Library        R                        �   �      n�         n�    �   ~   �?N �     �?N �   �   �   �  � ��-      � = Generic Library        T                        �   �   �?N �     �?N �   �   �  � ��)     � = Generic Library        N                        �   �   �?N 6�     �?N 6�   �   �  � ��)     � A Generic Library        N �                       �         ��         ��    �   }   �?N ��     �?N ��   �   �  �  } ��-      ��� M Generic Library        G �                       �   �      �         �    �   �   �?N .�     �?N .�   �   �  �  � ��;      � = Generic Library        J �                       �   �   �?N ��     �?N ��   �   �  � ��)     � ] Generic Library        I                        �         ^          ^     �   �   �?N       �?N     �   �  �   � ��M       � M Generic Library        E �                       �   �      �'         �'    �   �   �?N B�     �?N B�   �   �  �  � ��;      � = Generic Library        G                        �   �   �?N 
0     �?N 
0   �   �  � ��)     � = Generic Library        E                        �   �   �?N f�     �?N f�   �   �  � ��)     ��� M Generic Library       & 6 �                       �   �      �y         �y    �   �   �?N �}     �?N �}   �   �  �  � ��;      � M Generic Library       ! < �                       �   �      �l         �l    �   �   �?N q     �?N q   �   �  �  � ��;      � = Generic Library        A �                       �   �   �?N }     �?N }   �   �  � ��)     � A Generic Library        ?                        �   �      Z�         Z�    �   �   �?N 
�     �?N 
�   �   �  �  � ��-      � = Generic Library        <                        �   �   �?N �     �?N �   �   �  � ��)     � ] Generic Library        @                        �         �b         �b    �   �   �?N �^     �?N �^   �   �  �   � ��M       � A Generic Library        : �                       �   �      �|         �|    �   �   �?N �     �?N �   �   �  �  � ��-      � A Generic Library        9                        �         n�         n�    �   �   �?N �     �?N �   �   �  �   � ��-      � = Generic Library        7                        �   �   �?N       �?N     �   �   � ��)     � = Generic Library        5                        �   �   �?N 27     �?N 27   �   �  � ��)     � A Generic Library        5 �                       �   �      �         �    �   �   �?N &     �?N &   �   �  �  � ��-      � A Generic Library        4                        �   �      ��         ��    �   �   �?N ��     �?N ��   �   �  �  � ��-      � M Generic Library       ! 0                         �   �      �d         �d    �   �   �?N T�     �?N T�   �   ,  �  � ��;      ����� M Generic Library        �                        �         �         �    �   (   �?N ��     �?N ��   �   �   j  h ��;      � = Generic Library        �                        �   '   �?N �     �?N �   �   i  f ��)     � M Generic Library        j                         �         �         �    �   �   �?N      �?N    �   �  ]  � ��;      ��� M Generic Library       & ( �                       �   �      0h         0h    �   �   �?N <m     �?N <m   �   �  �  � ��;      � M Generic Library       ! % �                       �   �      *0         *0    �   �   �?N 65     �?N 65   �   �  �  � ��;      � = Generic Library        .                        �   �   �?N B9     �?N B9   �   �  � ��)     � A Generic Library        , �                       �   �      
[         
[    �   �   �?N >�     �?N >�   �   �  �  � ��-      � = Generic Library        , �                       �   �   �?N �u     �?N �u   �   �  � ��)     � ] Generic Library        +                        �         r�         r�    �   �   �?N ғ     �?N ғ   �   �  �   � ��M       � M Generic Library        '                        �         ��         ��    �   �   �?N n�     �?N n�   �   �  �  � ��;      � = Generic Library        k �                       �   z   �?N 
7     �?N 
7   �   �  � ��)     � = Generic Library        ( �                       �   �   �?N r     �?N r   �   �  �  ��)     � A Generic Library        " �                       �   �      �K         �K    �   �   �?N Ҵ     �?N Ҵ   �   �  �  � ��-      � = Generic Library        #                        �   �   �?N �     �?N �   �   �  � ��)     � M Generic Library        # �                       �                        �   �   �?N B�     �?N B�   �   �  �   � ��;      ��� = Generic Library        !                        �   �   �?N ��     �?N ��   �   �   ��)     � M Generic Library       &  �                       �   �      N         N    �   �   �?N �M     �?N �M   �   �  �  � ��;      � M Generic Library       !  �                       �   �      &�         &�    �   �   �?N ֎     �?N ֎   �   �  �    ��;      � M Generic Library       !  �                       �   �      ��         ��    �   �   �?N ��     �?N ��   �     �  � ��;      � = Generic Library                                �   �      ��         ��    �      ��)     � = Generic Library                                �   �   �?N bq     �?N bq   �   �    ��)     � = Generic Library                                �   �   �?N �     �?N �   �      ��)     � A Generic Library         �                       �         
�         
�    �   �   �?N ��     �?N ��   �        ��-      � A Generic Library         �                       �   �      X�         X�    �   �   �?N ��     �?N ��   �        ��-      � A Generic Library                                �         �         �    �   �   �?N \�     �?N \�   �   	  �    ��-      � A Generic Library         �                       �         h�         h�    �   �   �?N HT     �?N HT   �     
   ��-       A Generic Library         �                       �   �      �-         �-    �   �   �?N ~�     �?N ~�   �       � ��-      = Generic Library                                �   �   �?N ��     �?N ��   �      ��)     M Generic Library                                �   �      �#         �#    �   �   �?N v�     �?N v�   �         ��;      = Generic Library                                �   �   �?N �     �?N �   �   "  # ��)     � �    ��   �    �     ! ��     �    �   �    �    �    �    �   �    �    �    �    �    �    �    �    �    z    r    �    l    e    ]    K    G   v    ~    �    �    �    �    �     ! ��     �    �    �    �    �    �   �    �   �    �   �    �    �   �   �   �   r   l   h    e   \    X    Q    J    v   }    {    �   �    �    �    ! ��  �    �   �   �    �   �   �    �    �   �    �    �   �    �   �   �    �    �    �    s    m    [    Y   P    N    �    x    �    �    �   �   �    # ��     �   �    �    �    �    �    �    �   �    �   �   �    �   �   �   �    �   �   w    �   m   g    ]   \   W    Q   L   I    u   }   {   �   �      F    P      F   O      F    ��     G    H    	  G    M   
  H    J      H   I      K    L      L    M      M    O     N    O      P   Q      T    U      T   Y      T    ��  ��    U    ]      U   V      V    \      V   [      W    Z     X    Z      Y    Z      c    j      c   d      c    ��    d    i      d   f       e    f    !  f   g    "  h    i   #  i    m    $  j    n    %  j   k    &  k    l    '  n    �    (  n   �    )  p    t    *  p   q    +  p    ��  ,  q    r    -  q   s    .  t    x    /  t   u    0  u    v    1  w    x   2  z    |    3  {    |   4  |        5  }    ~   6  ~       7      �   8  �    ��  9  �    �    :  �   �    ;  �    ��  <  �    �    =  �   �    >  �    ��  ?  �    @  �   A  �   B  �   C  �    D  �    �    E  �    �   F  �    �    G  �   �    H  �    ��  I  �    �    J  �   �    K  �    �    L  �    �    M  �   �    N  �    �    O  �   �    P  �    �� 	 Q  �    �    R  �   �    S  �    �    T  �   �    U  �    �   V  �    �    W  �    �    X  �    �    Y  �    �    Z  �    �   [  �    �    \  �   �    ]  �    �    ^  �    �    _  �   �    `  �    �� 
 a  �    �    b  �   �    c  �    �   d  �    �    e  �    �    f  �   �    g  �    ��  h  �    �    i  �    �   j  �    �    k  �    �    l  �    �    m  �    �    n  �   �    o  �    ��  p  �    �    q  �   �    r  �    �    s  �    �    t  �   �    u  �    �    v  �    �    w  �    �    x  �   �    y  �    �    z  �   �    {  �    �   |  �    ��  }  �    �    ~  �   �      �    ��  �  �   �    �  �    �    �  �    �    �  �   �    �  �    ��  �  �    �    �  �    �    �  �   �    �  �    �    �  �   �    �  �    ��  �  �    �    �  �   �    �  �    �    �  �    �   �  �    �   �  �    �    �  �    �   �  �    �    �  �    �   �  �    �   �  �    �    �  �    �    �  �   �    �  �    ��  ��  �  �    �    �  �   �    �  �    �   �  �    �    �  �    �    �  �    �    �  �    �    �  �   �    �  �    �    �  �    �    �  �   �    �  �    ��  �  �    �    �  �   �    �  �        �  �   �    �  �    �   �  �    �    �  �    �    �  �    �    �         �        �         Generic Library         '        �         �    �        L-P                            Generic Library                  ��         ��    �   F     L-O                            Generic Library                 x�         x�    �   (     L-N                            Generic Library                 2�         2�    �        L-J                            Generic Library                  �         �    �   '     L-K                            Generic Library         '        �+         �+    �        L-L                            Generic Library         .        ��         ��    �        L-M                            Generic Library         .        V�         V�    �   Q     L-I                            Generic Library         '        ~         ~    �   T     L-H                            Generic Library                 f&         f&    �        L-F                            Generic Library                  �u         �u    �   +     L-G                                                                                                            	    	         
                       
                 	         
                                                                                      A (     ��   ����    # ! �� " ! ������������������������������������������ 
 N   P   % W !  X "  K #  L $ 1 [ % - Z & ) Y ' > V ( 9 U ) 8 S *   + "  ,   -    . 6 M / 4 R 0    1 5 O 2 T K 3 Q L 4 . M 5 + N 6 * O 7 ' P 8 & R 9  S :  U ;  V <  W = 	 X > F Y ?  Z @  [ \ A           0            -           ,           +           *   ��                .        @    '        ?   	        =   
                   "           #    .        !    '        <   ���������� .        ;    '        :             9       	                                                         ,          *     	                 0                            -   !  	        "       +   #  	          $    
           %  
          &          8   '          7   (               )      
  &   * '        6  
 +          5   ��-      	  %   . .        4  	 ����1        $   ����4        /   5        1  
 6        .  	 ��8        )   9        (   ��������>         '   ��������������F          >   ��������K '     2 "   L .     3 #   M .     4 .  	 N       5    O '     6 1  
 P   	    7    Q .        3   R       8 /   S       9 )   T '        2   U '     : (   V .     ; '   W ' 
    <     X .     ! =   Y       > &   Z '     ? %   [ .     @ $             A     B     C     D     E     L-Z     L-Y     L-X   	  L-V 	 	 
  L-R 
 
   L-S     L-T     L-U     L-Q  ��   L-P     L-O     L-N     L-J     L-K     L-L     L-M     L-I     L-H     L-F     L-G                                 	   
                            
   	                + V�      �An                                                         