 
 	    Generic Library                                   �          A0                            Generic Library                                  �        A1                            Generic Library                                  �        B0                            Generic Library                                  �        B1                            Generic Library                                  �    	    Ctrl0                         Generic Library         '        H8         H8    �        Z0                           ��  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   	  Generic Library         '        �r         �r    �        Z1                                                                                                 	      ��������                	   
                          	                                 
   ��                        ����         	    ��	           ��                                  �� '                 
                           '   	                                                	                                                                      ��       A0      A1     B0     B1     Ctrl0     Z0   	  Z1 	                           L ��       �An                                                         