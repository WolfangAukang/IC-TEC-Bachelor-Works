 q i    Generic Library                                   �         A                             Generic Library          
                        �        D                             Generic Library                                  �   	     B                             Generic Library                                  �   )     C                            M Generic Library       &                          �         N�         N�    �         ��         ��    �      *     ��;        Generic Library         . E 4      ��         ��    �        W                              Generic Library         . 1 &      p         p    �        U                             M Generic Library       & 	                        �         V�         V�    �         Ʒ         Ʒ    �   :   4     ��;        Generic Library         1  
      �E         �E    �        T                            	 M Generic Library       +                         �   	      ��         ��    �   
      ~�         ~�    �           ��;      
 M Generic Library       &                         �         *�         *�    �   	      ��         ��    �   K   R     ��;       M Generic Library       +                         �                      �         �         �    �            ��;       M Generic Library       &                          �         $�         $�    �         �         �    �   =   G     ��;        Generic Library         0        V�         V�    �        S                              Generic Library         ( X >      ��         ��    �   �     X                              Generic Library         - � a      >         >    �      	  Z                              Generic Library         - n M      �G         �G    �   
   
  Y                             = Generic Library                                �         �d         �d    �        ��)      = Generic Library                                �         $         $    �   +   ,  ��)      A Generic Library        
                        �         �         �    �         H          H     �   7      <  ��-       A Generic Library                                �         .�         .�    �         �&         �&    �      ,   3  ��-       = Generic Library                                �         �d         �d    �   B   "  ��)      = Generic Library                                �         $         $    �   E     ��)      = Generic Library                                �         $         $    �         ��)      A Generic Library                                �         X^         X^    �         ��         ��    �      H   C  ��-       A Generic Library                                �         ��         ��    �         Z�         Z�    �   "      D  ��-       A Generic Library        !                        �         ��         ��    �         Q         Q    �   L   O   P  ��-       = Generic Library        !                        �         2E         2E    �   N   L  ��)      D Generic Library        &                        �         �&         �&    �         H          H     �         (         (    �   U   e   T   �  ��0       D Generic Library        *                        �         ��         ��    �         4�         4�    �         ��         ��    �   {   V   |     ��0       D Generic Library        .                         �         ��         ��    �         �          �     �         |          |     �   }   ~   [   ]  ��0       A Generic Library        2                        �         (�         (�    �         ,�         ,�    �   d   c   b  ��-        A Generic Library        6                         �   !      ��         ��    �   "      X�         X�    �   a   `   �  ��-      ! = Generic Library        &                         �         �         �    �   j   m  ��)     " = Generic Library        '                        �         nn         nn    �   k   g  ��)     # = Generic Library        (                        �         Ve         Ve    �   l   i  ��)     $ = Generic Library        *                         �         �$         �$    �   o   n  ��)     % = Generic Library        /                        �                      �   r   q  ��)     & = Generic Library        2                        �         �         �    �      �  ��)     ' = Generic Library        4                        �         @�         @�    �   �   t  ��)     ( = Generic Library        6                        �          ��         ��    �   v   �  ��)     ) = Generic Library        8                        �   !      H�         H�    �   �   x  ��)     * M Generic Library        (                        �         �U         �U    �   #      XU         XU    �   z   �   Y  ��;      + M Generic Library        0                        �         �F         �F    �   $      hF         hF    �   �   �   �  ��;      , M Generic Library       $ , #                       �   $      9         9    �   %      �8         �8    �   �   �   �  ��;      - M Generic Library       ) 0 %                       �   "      �         �    �   &      ��         ��    �   �   �     ��;      . D Generic Library        ; '                       �         �&         �&    �   (      H          H     �   )      (         (    �   �   �   �   �  ��0      / D Generic Library        ?                        �   *      ��         ��    �         4�         4�    �   +      ��         ��    �   �   �   �   �  ��0      ��1 A Generic Library        G ,                       �         (�         (�    �   -      ,�         ,�    �   �   �   �  ��-      2 A Generic Library        K                         �         ��         ��    �   .      X�         X�    �   �   �   �  ��-      3 = Generic Library        ;                         �   '      H�         H�    �   �   �  ��)     4 = Generic Library        =                        �   (      H�         H�    �   �   �  ��)     5 = Generic Library        @                        �   *      H�         H�    �   �   �  ��)     6 = Generic Library        E                        �   /      H�         H�    �   !  �  ��)     7 = Generic Library        G                        �   ,      H�         H�    �   �   �  ��)     8 M Generic Library        = )                       �   +      �         �    �   0      (�         (�    �   �   �   �  ��;      ��: M Generic Library        E 1                       �   -      �j         �j    �   2      �j         �j    �   �   �   �  ��;      ; M Generic Library       $ A 0                       �   2      �         �    �   3      l         l    �   �   �   �  ��;      < M Generic Library       ) D 3                       �   .      |         |    �   4      ��         ��    �   �   �     ��;      = A Generic Library        Q 5                       �   6      ��         ��    �   7      p�         p�    �   �   �   �  ��-      > A Generic Library        U 8                       �         ��         ��    �   9      z�         z�    �   �   �   �  ��-      ? A Generic Library        Y                         �         \�         \�    �   :      �         �    �   �   �   �  ��-      @ A Generic Library        ]                         �         ��         ��    �   ;      Z�         Z�    �   �   �   �  ��-      A = Generic Library        Q                        �   5      H�         H�    �   �   �  ��)     B = Generic Library        S                        �   6      �B         �B    �   �   �  ��)     C = Generic Library        U                        �   8      ��         ��    �   �   �  ��)     ��E M Generic Library        S 7                       �   9      L         L    �   <      NC         NC    �   �   �   �  ��;      F M Generic Library        [ :                       �   ;                   �   =      �         �    �   �   �   �  ��;      G M Generic Library       # W <                       �   =      ��         ��    �   >      >�         >�    �   �   �   �  ��;      ������K A Generic Library        n ?                       �         (�         (�    �   @      ,�         ,�    �   �   �   �  ��-      L A Generic Library        r                         �   A      ��         ��    �   B      X�         X�    �   �   �    ��-      ����O = Generic Library        t                        �   A      �[         �[    �   �   �  ��)     P = Generic Library        n                         �   ?      �         �    �     �  ��)     Q A Generic Library        b C                       �   D      �_         �_    �   E      �         �    �       �  ��-      R = Generic Library        j                        �   F      *{         *{    �       ��)     S = Generic Library        f                        �   G      f#         f#    �     	 ��)     T = Generic Library        d                        �   D      �8         �8    �      ��)     U = Generic Library        b                        �   C      �         �    �      ��)     V M Generic Library        d E                       �   H      X�         X�    �   I      �$         �$    �        ��;      W M Generic Library        l J                       �   @      J'         J'    �   K      �&         �&    �        ��;      X M Generic Library       # h I                       �   K      Fo         Fo    �   L      �n         �n    �        ��;      Y M Generic Library       ( m L                       �   B      �a         �a    �   M      Da         Da    �       
  ��;      Z D Generic Library        w N                       �   O      P         P    �   P                     �   Q      �         �    �          D ��0      [ A Generic Library        f G                       �         ^I         ^I    �   H      �         �    �   	    �  ��-      \ D Generic Library        { R                       �         R�         R�    �         m         m    �   S      �%         �%    �   %  R  S    ��0      ] D Generic Library         T                       �         N          N     �   U      FS         FS    �   V      p�         p�    �   &   U  +  ( ��0      ^ D Generic Library        �                        �   W      j�         j�    �         �         �    �   X      ��         ��    �   W  .  Y  , ��0      _ D Generic Library        �                         �         ��         ��    �   Y      �I         �I    �   Z      �         �    �   Z  [  "  1 ��0      ` A Generic Library        �                         �   [      u         u    �   \      l�         l�    �   ]     7 ��-      a = Generic Library                                 �   T      �         �    �   T  &  ��)     b = Generic Library        {                        �   R      &�         &�    �   Q  % ��)     c = Generic Library        y                        �   P      �=         �=    �   P   ��)     d = Generic Library        x                        �   O      &}         &}    �   <   ��)     e = Generic Library        w                        �   N      R         R    �   M    ��)     f = Generic Library        �                        �   U      b�         b�    �   V  + ��)     g = Generic Library        �                        �   W      �         �    �   X  . ��)     h = Generic Library        �                        �   [      �         �    �       ��)     i A Generic Library        j F                       �         ��         ��    �   J      n�         n�    �     �   �  ��-      j A Generic Library        C                         �   /      Z�         Z�    �   1      *         *    �   �   $  �  ��-      k = Generic Library        �                        �   Y      H          H     �   \  " ��)     l M Generic Library        y Q                       �   S      �         �    �   ]      ��         ��    �   2  @  N ��;      m M Generic Library        � V                       �   X      �H         �H    �   ^      �B         �B    �   B  C  A ��;      n M Generic Library        � Z                       �   \      vp         vp    �   _      ��         ��    �   0  E  O ��;      o M Generic Library       # } ]                       �   ^      ��         ��    �   `      l�         l�    �   H  I  J ��;      p M Generic Library       ( � `                       �   _      
"         
"    �   a      FS         FS    �   F  K    ��;      b b             $        3    j    2    ?    @    P    a    _    `    L    !                      #          )    4    /   B    C    [   c    \   f    ^   k    i                      &    (    .   /    7    A    @   U    S    K   e    b    ^    _   O    6                          %    '    5    1   2   >   ?   T    R    d    \   ]   g    h       "                                               	        	  	   
    
  	          
          
                                                                                          !         "         #          *          $          *        %          +          &         '          +           (    !      )    "       -   #  *    ,    $  +    ,   %  ,    -    &  -        '  .    3    (  .   4    )  .    8    *  /   5    +  /    8   ,  1    7    -  1    :   .  2    <   /  6    j   0  8    ;    1  :    j    2  :    ;   3  ;    <    4  <        5  =    A    6  =   B    7  =    E    8  >    C    9  >    E   :  ?    F    ;  @    F   <  E    G    =  F    G   >  G        ?  K    P    @  K    W   A  L   O    B  L    Y   C  Q    U    D  Q   T    E  Q    V    F  R    i    G  S    [    H  V   [    I  V    X    J  W    i    K  W    X   L  X    Y    M  Y        N  Z    e    O  Z   d    P  Z   c    Q  Z    l    R  \    b    S  \    l   T  ]    a    U  ]   f    V  ]    m    W  ^   g    X  ^    m   Y  _   k    Z  _    n    [  `   h    \  `    n   ]  l    o    ^  m    o   _  n    p   `  o    p    a  p        � �   .   1 4  1 3  / .  / 6 �� ! *  2 B  #  	 - + 
 � � �� 	   ( 2  %    A  � �   #  # 9  9 =      @ ��       5 0  % 5   %   /  6 7  8   5 -   0 8 !   "   # ( > $ ; : % ; < & ) ( ' ! > (  E )  M * F D + 2 ? , ?   - � � . A H / J K 0 J C 1 F G 2 M N 3 A I 4 I O 5 @ R 6 P Q 7 @ Q 8 9 ^ ��: ? f ��< M h = h l ����@ i T A ^ S B S o C f W D p r E n { F p W G W V H h X I X | J S Z K Z } L q ~ M X \ N \ [ O I s P s  Q p u R u � S � d T t c U s w V w v W \ y X y � Y � a Z x ` [ � z \ �  ] Y � ^ ] � _ � b ` � � a � _ b � � c � _ d Z � e � � f � � g y � h � � i � � j w � k � � ��m � � n u � o � � p � !q � � r � � s � � t � � u g e v � � w � � x � � y � $z D2{ � � | � � } � � ~ � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � #� � � � � � � � � � � � � � f k � m U � ^ j � � � IA� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � NH� 
� � � � ;� � � �  � ;&� � � � � � � 
� 
� � � � � � G� � � � � � � � � � :� 8� � G9� 84� :'� � � � � � � � � � � � � � � � � � (B� C,� 10� E7� JF� KL� OL� ^� GM� � ^� ;<� ' ?� :P� � � � 9Q� � � � &R� � � � 'S� 65� 8T� &*� *U� ')� )V� 9-� -W� *=� =X� )/� /Y� � � � 4Z� >3� 3[� /?� ?\� 45� 5]� =^� -3_J  + 
          +                                           +                       +            	            &            	 	           
 - o      Y       M               0 	               - �      p       a  	               x  Z    e       N ����       ( )     �  `   h       [            �� . F      <       4  . 2      -       &  +        "    1        !  
  +   	      	  +   	     "    0   	     !  
   ,       \                    +   
       	           ,   ! #      '   "                #            ��%           &  �  a    ]       T '  �    �   (  	     & #   ) 	 	       &   * &          +         	   ,               -       	   .           /           0           1 $         2        +   3 $           4 &          5           6          7            8           9        8    : & 
       $   ; ! 
    $ %   < !        %   = &            > # 	    ' #   ?      + , :   @       7 5   A       . 3   B            C         0   D         *   E         (   F      1 *   G &       1   H        .   I  $    3 4 O   J      / 0   K &   
     /   L  "              M  "    ) 2 <   N  "       2   O  $      4   P  #       6   Q   #    6 7   R &   
    5   S  +    A B J    T  )      @   U  '       �   V  ,      G   W  ,    F C G   X  -    H I M   Y $ *  *     ]  # Z  /    J K d    [  1      N   \  1    M N W   ]  0       ^   ^  '    8 A �    _ ) 8    a c  " `  9       Z  ! a  7        Y    b  4       _   c  5      T   d  3       S   e  (      u   f  (    : C �   g  (  "     u   h  )    < = H   i  )  #     @   j  '  !     �    k  (  "     �   l  )  #     =   m  '  !     �   n  +  $     E   o  +  $     B    p  0    D F Q   q  0  %     L   r  0  %     D   s  3    O P U   t  5  '     T   u  5    Q R n   v  7  (     V   w  7    U V j   x  9  )     Z  ! y  9    W X g   z  )  *     [   {  +       E   |  -      I   }  /       K    ~  0      L     3  &     P   �  5  '     R   �  3  &     S   �  9  )     X   �  7  (     Y    �  +  *    \   �  1  +     ^   �  3  +    _   � $ 2  +     `  $ �  8        a  " � $ -  ,     ]  # � $ /  ,    `  $ � ) 3  -    c  " �  (       [   � ) 1  -     b  % �  =    j k �   �  <  .     f  ' � ) .  ,     b  % �  >  .    i  ( �  =  .     �  ) �  @    m � r   �  A  /    x  * �  B    q � �   �  A  /     �  + �  D    v w �    �����  E  j     �  1 �  H  1     |  , �  J    } ~ �   �  I  1     �  - �  L    � � �    �  N    � � �   � ) M    � �  . �  >  4     h   �  <    d e v    �  >    g h �   �  =  .    k   �  A    n o }   �  F  6     � y  / ���  H  7     {   �  H    { s �   �  J  1    ~   �  <  3     e    �  <  3     f  ' �  >  4     i  ( �  @  /     m   �  A  5     o   �  B  /    q   �����  D  j     w    �  A  5     x  * �  H  7     |  , �  L  2     �    �  N  2    �   �  @  8    �  + �  F  :     �  1 � $ D  ;    �  2 �����  F    r s p   �  H  :    �  - � $ B  ;     �  0 � $ G  :     �  2 �  >  8     �  ) � ) E  <     �  3 �  M  2     �  . � $ ?  8     �  0 �  T  =   B       6 �  R    - � �   � ) C  ;     �  3 � ) G  <    �  . �  [  ?     �  : �  V  C    >       8 ���  S  =     �  7 �  `  @    
   �  ^  @         �  _  @     �  ; �  \    t � �   �  Z  ?         � # X  G     �  < �  R  =    A       5 �  T    � � �   �  X  >    �   �  V  C     �   �  R  A     -   �  T  B     �   �  V    � � �   �  X    � � �   �  Z    �  �    �  \  ?    t   �  ^     � �    �  `    
 � �   �  T  E     �  7 �  V  E    �  9 � # ]  F     �  = �  \  F     �  : �  ^  F    �  ; � ( Y      G       > �  W  >     �  9 � # Z  G    �  = �  �    �   � # U  E     �  < �������  d  Q     �  E �������  h  [     �  H �������  l  i     �  J �  o  K    P       ? �  u  O     �   �  p  K     �  @ �  s    � � �    �  u  L   O       A � ( t    � �  B �  s  L     �    �  q    � � �   �  q  K    �   �  o    � � �    �  m  i    �     k  R     �    i  [    �    g  S     �    e  Q   T       D  c  Q    U       C  e  T     �    c  U     �    u    � � �    k  R    i       F 	 g  S    [       G 
 g    � � �    e    � � �    c    � � �    i    � � �    k    � � �    m    � � �    o  P     �     m  W     �  J  e  V     �  E # f  V     �  I  o  W    �  @ # k  X    �  K # n  W     �  K ( n  Y     �  L # i  X     �  I ( j  X     �  L  t  L     �  B  �  h     �    g  V    �  H ( p  Y    �  B  y  Z   d       O  z  Z   c       P   }  \       S ! F  6     p   " �  k    _      Y # F    �  / $ F  j    y  / % |  \    b       R & }    � � �   ' ~    � � �   ( �  ]     �  V ) �    � � �   * �    � � �   + �  ]   f       U , �  ^     �  X - �    � � �   . �  ^   g       W / �    � � �   0 �  n     �  Z 1 �  _     �  Z 2 z  l     z  Q 3 �    � � �   4 �    � � �    5 �    � � �    6 �    �    7 �  `     �  \ 8 �    � � �    9 |    � � �   : z    � � �   ; y    � � �   < y  d     �   = �    � � �   > �    �   ? �    � � �   @ |  l      S A# �  m     �  ^ B �  m     �  V C �  m    �  X D y  Z     z  Q E �  n    �  \ F( �  p     �  ` G x    � � �   H# ~  o     �  ] I# �  o    �  ^ J(   o     �  ` K( �  p    �  _ L( �    � �  _ M x  e     �   N# {  l     �  ] O# �  n     �  _ P z  c     �   Q |  b     �   R }  \    �   S ~  \    �   T �  a     �    U �  ]    �   V �  f     �   W �  ^     �   X �  g     �   Y �  ^    �   Z �  _     �    [ �  _    �   \ �  k     �   ] �  `     �    ^ �    � � �     �� )  =  
 201308685  )  =  q Kafay Rafael Ng Zhao          2013102458                     Fundamentos de Organizaci�n de Computadores Grupo 2  )  =   7 Segmentos        A      D     B     C     S     T     U     W     X  	   Z  
   Y                                 	 	  
 
   J N�       �An                                                         