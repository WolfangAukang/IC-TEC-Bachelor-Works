      Generic Library                               �         ��         ��    �         ��         ��    �         ��         ��    �         �         �    �         ě         ě    �         �         �    �         ��         ��    �         ��         ��    �   	       8          8    �   
      �f         �f    �                              ��  @cQ 086585S.CKT& C:\USERS\LEEECHER\DOCUME~1\086585S.CKT 086585S.CKTA �p W�    D �p W�   B �p W�   C �p W�   W �p W�    U �p W�   T �p W�   S �p W�   X �p W�   Z �p W�   Y �p W�   ����������������������  �� �� �� ��4 ��& ��
 �� ��> ��a ��M ��q ^ �������� M Generic Library       &                          �         N�         N�    �         ��         ��    �      *     ��;      ���� M Generic Library       & 	                        �         V�         V�    �         Ʒ         Ʒ    �   :   4     ��;      ��	 M Generic Library       +                         �   	      ��         ��    �   
      ~�         ~�    �           ��;      
 M Generic Library       &                         �         *�         *�    �   	      ��         ��    �   K   R     ��;       M Generic Library       +                         �                      �         �         �    �            ��;       M Generic Library       &                          �         $�         $�    �         �         �    �   =   G     ��;      �������� = Generic Library                                �         �d         �d    �        ��)      = Generic Library                                �         $         $    �   +   ,  ��)      A Generic Library        
                        �         �         �    �         H          H     �   7      <  ��-       A Generic Library                                �         .�         .�    �         �&         �&    �      ,   3  ��-       = Generic Library                                �         �d         �d    �   B   "  ��)      = Generic Library                                �         $         $    �   E     ��)      = Generic Library                                �         $         $    �         ��)      A Generic Library                                �         X^         X^    �         ��         ��    �      H   C  ��-       A Generic Library                                �         ��         ��    �         Z�         Z�    �   "      D  ��-       A Generic Library        !                        �         ��         ��    �         Q         Q    �   L   O   P  ��-       = Generic Library        !                        �         2E         2E    �   N   L  ��)      D Generic Library        &                        �         �&         �&    �         H          H     �         (         (    �   U   e   T   �  ��0       D Generic Library        *                        �         ��         ��    �         4�         4�    �         ��         ��    �   {   V   |     ��0       D Generic Library        .                         �         ��         ��    �         �          �     �         |          |     �   }   ~   [   ]  ��0       A Generic Library        2                        �         (�         (�    �         ,�         ,�    �   d   c   b  ��-        A Generic Library        6                         �   !      ��         ��    �   "      X�         X�    �   a   `   �  ��-      ! = Generic Library        &                         �         �         �    �   j   m  ��)     " = Generic Library        '                        �         nn         nn    �   k   g  ��)     # = Generic Library        (                        �         Ve         Ve    �   l   i  ��)     $ = Generic Library        *                         �         �$         �$    �   o   n  ��)     % = Generic Library        /                        �                      �   r   q  ��)     & = Generic Library        2                        �         �         �    �      �  ��)     ' = Generic Library        4                        �         @�         @�    �   �   t  ��)     ( = Generic Library        6                        �          ��         ��    �   v   �  ��)     ) = Generic Library        8                        �   !      H�         H�    �   �   x  ��)     * M Generic Library        (                        �         �U         �U    �   #      XU         XU    �   z   �   Y  ��;      + M Generic Library        0                        �         �F         �F    �   $      hF         hF    �   �   �   �  ��;      , M Generic Library       $ , #                       �   $      9         9    �   %      �8         �8    �   �   �   �  ��;      - M Generic Library       ) 0 %                       �   "      �         �    �   &      ��         ��    �   �   �     ��;      . D Generic Library        ; '                       �         �&         �&    �   (      H          H     �   )      (         (    �   �   �   �   �  ��0      / D Generic Library        ?                        �   *      ��         ��    �         4�         4�    �   +      ��         ��    �   �   �   �   �  ��0      ��1 A Generic Library        G ,                       �         (�         (�    �   -      ,�         ,�    �   �   �   �  ��-      2 A Generic Library        K                         �         ��         ��    �   .      X�         X�    �   �   �   �  ��-      3 = Generic Library        ;                         �   '      H�         H�    �   �   �  ��)     4 = Generic Library        =                        �   (      H�         H�    �   �   �  ��)     5 = Generic Library        @                        �   *      H�         H�    �   �   �  ��)     6 = Generic Library        E                        �   /      H�         H�    �   !  �  ��)     7 = Generic Library        G                        �   ,      H�         H�    �   �   �  ��)     8 M Generic Library        = )                       �   +      �         �    �   0      (�         (�    �   �   �   �  ��;      ��: M Generic Library        E 1                       �   -      �j         �j    �   2      �j         �j    �   �   �   �  ��;      ; M Generic Library       $ A 0                       �   2      �         �    �   3      l         l    �   �   �   �  ��;      < M Generic Library       ) D 3                       �   .      |         |    �   4      ��         ��    �   �   �     ��;      = A Generic Library        Q 5                       �   6      ��         ��    �   7      p�         p�    �   �   �   �  ��-      > A Generic Library        U 8                       �         ��         ��    �   9      z�         z�    �   �   �   �  ��-      ? A Generic Library        Y                         �         \�         \�    �   :      �         �    �   �   �   �  ��-      @ A Generic Library        ]                         �         ��         ��    �   ;      Z�         Z�    �   �   �   �  ��-      A = Generic Library        Q                        �   5      H�         H�    �   �   �  ��)     B = Generic Library        S                        �   6      �B         �B    �   �   �  ��)     C = Generic Library        U                        �   8      ��         ��    �   �   �  ��)     ��E M Generic Library        S 7                       �   9      L         L    �   <      NC         NC    �   �   �   �  ��;      F M Generic Library        [ :                       �   ;                   �   =      �         �    �   �   �   �  ��;      G M Generic Library       # W <                       �   =      ��         ��    �   >      >�         >�    �   �   �   �  ��;      ������K A Generic Library        n ?                       �         (�         (�    �   @      ,�         ,�    �   �   �   �  ��-      L A Generic Library        r                         �   A      ��         ��    �   B      X�         X�    �   �   �    ��-      ����O = Generic Library        t                        �   A      �[         �[    �   �   �  ��)     P = Generic Library        n                         �   ?      �         �    �     �  ��)     Q A Generic Library        b C                       �   D      �_         �_    �   E      �         �    �       �  ��-      R = Generic Library        j                        �   F      *{         *{    �       ��)     S = Generic Library        f                        �   G      f#         f#    �     	 ��)     T = Generic Library        d                        �   D      �8         �8    �      ��)     U = Generic Library        b                        �   C      �         �    �      ��)     V M Generic Library        d E                       �   H      X�         X�    �   I      �$         �$    �        ��;      W M Generic Library        l J                       �   @      J'         J'    �   K      �&         �&    �        ��;      X M Generic Library       # h I                       �   K      Fo         Fo    �   L      �n         �n    �        ��;      Y M Generic Library       ( m L                       �   B      �a         �a    �   M      Da         Da    �       
  ��;      Z D Generic Library        w N                       �   O      P         P    �   P                     �   Q      �         �    �          D ��0      [ A Generic Library        f G                       �         ^I         ^I    �   H      �         �    �   	    �  ��-      \ D Generic Library        { R                       �         R�         R�    �         m         m    �   S      �%         �%    �   %  R  S    ��0      ] D Generic Library         T                       �         N          N     �   U      FS         FS    �   V      p�         p�    �   &   U  +  ( ��0      ^ D Generic Library        �                        �   W      j�         j�    �         �         �    �   X      ��         ��    �   W  .  Y  , ��0      _ D Generic Library        �                         �         ��         ��    �   Y      �I         �I    �   Z      �         �    �   Z  [  "  1 ��0      ` A Generic Library        �                         �   [      u         u    �   \      l�         l�    �   ]     7 ��-      a = Generic Library                                 �   T      �         �    �   T  &  ��)     b = Generic Library        {                        �   R      &�         &�    �   Q  % ��)     c = Generic Library        y                        �   P      �=         �=    �   P   ��)     d = Generic Library        x                        �   O      &}         &}    �   <   ��)     e = Generic Library        w                        �   N      R         R    �   M    ��)     f = Generic Library        �                        �   U      b�         b�    �   V  + ��)     g = Generic Library        �                        �   W      �         �    �   X  . ��)     h = Generic Library        �                        �   [      �         �    �       ��)     i A Generic Library        j F                       �         ��         ��    �   J      n�         n�    �     �   �  ��-      j A Generic Library        C                         �   /      Z�         Z�    �   1      *         *    �   �   $  �  ��-      k = Generic Library        �                        �   Y      H          H     �   \  " ��)     l M Generic Library        y Q                       �   S      �         �    �   ]      ��         ��    �   2  @  N ��;      m M Generic Library        � V                       �   X      �H         �H    �   ^      �B         �B    �   B  C  A ��;      n M Generic Library        � Z                       �   \      vp         vp    �   _      ��         ��    �   0  E  O ��;      o M Generic Library       # } ]                       �   ^      ��         ��    �   `      l�         l�    �   H  I  J ��;      p M Generic Library       ( � `                       �   _      
"         
"    �   a      FS         FS    �   F  K    ��;      b b    ��       !    $        3    j    2    ?    @    P    a    _    `    L          ��          #          )    4    /   B    C    [   c    \   f    ^   k    i            ��        &    (    .   /    7    A    @   U    S    K   e    b    ^    _   O    6              ��          "    %    '    5    1   2   >   ?   T    R    d    \   ]   g    h                                                  	        	  	   
    
  	    ��    
          
             ��                                                                           !         "         #          *          $          *        %          +          &         '          +           (    !      )    "       -   #  *    ,    $  +    ,   %  ,    -    &  -    ��  '  .    3    (  .   4    )  .    8    *  /   5    +  /    8   ,  1    7    -  1    :   .  2    <   /  6    j   0  8    ;    1  :    j    2  :    ;   3  ;    <    4  <    ��   5  =    A    6  =   B    7  =    E    8  >    C    9  >    E   :  ?    F    ;  @    F   <  E    G    =  F    G   >  G    ��  ?  K    P    @  K    W   A  L   O    B  L    Y   C  Q    U    D  Q   T    E  Q    V    F  R    i    G  S    [    H  V   [    I  V    X    J  W    i    K  W    X   L  X    Y    M  Y    ��  N  Z    e    O  Z   d    P  Z   c    Q  Z    l    R  \    b    S  \    l   T  ]    a    U  ]   f    V  ]    m    W  ^   g    X  ^    m   Y  _   k    Z  _    n    [  `   h    \  `    n   ]  l    o    ^  m    o   _  n    p   `  o    p    a  p    ��    Generic Library                                   �         In0                           Generic Library                                  �        In1                           Generic Library                                  �        In2                           Generic Library          	                        �        In3                          s Generic Library                                   �         ��         ��    �   
      {         {    �   	      �         �    �         J�         J�    �         ��         ��    �         Z�         Z�    �                     
   ��                                                                                            	         
                         ��           
 	   
                               
                                      	 ��         	   ��   	         ��
                                                    
                                                	    
           	          ��         	            
                  
         
            
         � Pedro Henrique Rodriguez de Oliveira 2013086585 Fundamentos de Organizaci�n de computadoras Grupo 1 Encapsulado del 7 segmentos       In0     In1     In2     In3                   / R�       �An                                                         