      Generic Library                                   �         A                             Generic Library                                  �        B                             Generic Library                                  �        C                             Generic Library         &  	                       �        Y                              Generic Library         +                         �        X                             = Generic Library                                �      �?N ��     �?N ��   �   	     ��)      A Generic Library                                �         �         �    �      �?N B�     �?N B�   �         !  ��-       = Generic Library                                 �      �?N ��     �?N ��   �      
  ��)      = Generic Library        
                        �      �?N ��     �?N ��   �        ��)     	 ] Generic Library                                �         d�         d�    �      �?N �     �?N �   �           ��M       
 A Generic Library        	                        �          �         �    �      �?N B�     �?N B�   �            ��-       M Generic Library       !                         �         ,k         ,k    �   	   �?N �j     �?N �j   �            ��;       ] Generic Library                                �          d�         d�    �   
   �?N �     �?N �   �         "  ��M        = Generic Library         
                       �      �?N ��     �?N ��   �   "   '  ��)      A Generic Library                                 �         �         �    �      �?N B�     �?N B�   �   ,   '   +  ��-       M Generic Library       &                         �         ,k         ,k    �      �?N �j     �?N �j   �   )   -     ��;       A Generic Library                                 �         �         �    �      �?N B�     �?N B�   �   /   2   1  ��-                       
             	                  	                                                   	    
      
       	          
                                                $ $          	      *               	   
                $ #     (   0      !    0  * $      &      *  &   0 (  # ,  + )  . -   . 1 ! 
 2 "  % # % / 4 3      
          
                     &              	  +                             	                   
              	            
         !                 	  	          	                                                                  	                        	                     
  "       	         
  	    
          
                    !            !          !   
                                 !          !            "               
 #           $          %      " #   &          '                (           ) &           *  	         + %           ,             - &          . %          /          #   0            1 %            2         !   ��           A      B     C     Y     X                     & 5 �f      �An                                                          