      Generic Library                �j         �j    �         ��         ��    �         ��         ��    �         ��         ��    �         �         �    �      	   
       ��  �z[Q
 ALARMA.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\ALARMA.CKT
 ALARMA.CKTA �m W�    B �m W�   C �m W�   Y �m W�    X �m W�   ����������  �� �� ��	 �� ��  ���������� = Generic Library                                �      �?N ��     �?N ��   �   	     ��)      A Generic Library                                �         �         �    �      �?N B�     �?N B�   �         !  ��-       = Generic Library                                 �      �?N ��     �?N ��   �      
  ��)      = Generic Library        
                        �      �?N ��     �?N ��   �        ��)     	 ] Generic Library                                �         d�         d�    �      �?N �     �?N �   �           ��M       
 A Generic Library        	                        �          �         �    �      �?N B�     �?N B�   �            ��-       M Generic Library       !                         �         ,k         ,k    �   	   �?N �j     �?N �j   �            ��;       ] Generic Library                                �          d�         d�    �   
   �?N �     �?N �   �         "  ��M        = Generic Library         
                       �      �?N ��     �?N ��   �   "   '  ��)      A Generic Library                                 �         �         �    �      �?N B�     �?N B�   �   ,   '   +  ��-       M Generic Library       &                         �         ,k         ,k    �      �?N �j     �?N �j   �   )   -     ��;       A Generic Library                                 �         �         �    �      �?N B�     �?N B�   �   /   2   1  ��-           ��          
     ��      	          ��      	                                                   	    
      
       	      ��   
                                            ��    Generic Library                 ��         ��    �         "�         "�    �          ��         ��    �    
     Suceso                       ` Generic Library              4         4    �         �!         �!    �          �         �    �         $*         $*    �         �%         �%    �          �2         �2    �             ��	                                     Generic Library                                  �         TH         TH    �        Bips                          ` Generic Library               �         �    �         d;         d;    �         �?         �?    �         "�         "�    �           ��                                                                                          	   
         	                                                                                                 ��  	            	            
            ��                                    Suceso     Bips            ) 8 �i       �?N                                                          