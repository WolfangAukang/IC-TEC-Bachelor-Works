 �    Generic Library                                   �        A                             Generic Library                                  �   	     B                             Generic Library                                  �   )     C                             Generic Library          
                        �   �     D                             Generic Library                                  �       E                           ��������������������������������������������������������������������������������������������������������������������������������E  Generic Library         0       8         8    �   �     L-Z                          F M Generic Library       +                        �         �#         �#    �      �?N �     �?N �   �     �   �  ��;      G A Generic Library                               �         �[         �[    �   	   �?N Dj     �?N Dj   �   �   �   �  ��-      H A Generic Library        
                         �         X         X    �      �?N ��     �?N ��   �   �   �   �  ��-      I = Generic Library                               �      �?N ��     �?N ��   �   �   �  ��)     J = Generic Library                                 �   
   �?N J�     �?N J�   �     �  ��)     K = Generic Library        
                       �      �?N >     �?N >   �      ��)     L A Generic Library        
                       �         ��         ��    �      �?N >     �?N >   �        ��-      M M Generic Library       !                        �   	      ��         ��    �      �?N �C     �?N �C   �     �   �  ��;      N = Generic Library                               �      �?N B/     �?N B/   �   ^  	 ��)     O A Generic Library       & 
                       �         �o         �o    �      �?N �     �?N �   �     �    ��-      P A Generic Library                               �         �         �    �      �?N ��     �?N ��   �        ��-      Q ] Generic Library                               �         &1         &1    �      �?N �\     �?N �\   �        ��M       R  Generic Library         & �       ��         ��    �       L-Y                          S  Generic Library         & �       �         �    �       L-X                          T M Generic Library       ! �                        �         N�         N�    �      �?N �f     �?N �f   �         ��;      U M Generic Library        �                        �         V.         V.    �      �?N ޜ     �?N ޜ   �   #  !  " ��;      V A Generic Library        �                        �         �         �    �      �?N p.     �?N p.   �   $  4   ��-      W = Generic Library                                �      �?N &U     �?N &U   �   &  ' ��)     X = Generic Library        �                        �      �?N *     �?N *   �   -  ( ��)     Y A Generic Library        �                        �          �          �    �      �?N n�     �?N n�   �   +    ) ��-      Z A Generic Library        �                        �         �%         �%    �      �?N f!     �?N f!   �   (  '  + ��-      [ = Generic Library        �                        �      �?N v�     �?N v�   �     0 ��)     \ ] Generic Library        �                        �         ��         ��    �      �?N ��     �?N ��   �   3  2  $ ��M       ] A Generic Library        �                        �         ��         ��    �      �?N >�     �?N >�   �   <  8   ��-      ^  Generic Library         & �       8�         8�    �   9    L-V                          ��������c M Generic Library       ! �                        �         �r         �r    �      �?N �W     �?N �W   �   H  \  9 ��;      d M Generic Library        �                        �         ��         ��    �      �?N ��     �?N ��   �   I  Y  G ��;      e A Generic Library        �                        �         �1         �1    �       �?N N�     �?N N�   �   L  K  O ��-      f A Generic Library        �                         �   !      �W         �W    �      �?N F�     �?N F�   �   T  S  R ��-      g = Generic Library        �                        �   !   �?N ʎ     �?N ʎ   �   J  S ��)     h = Generic Library        �                        �   "   �?N ʎ     �?N ʎ   �   M  V ��)     i A Generic Library        � #                       �   "      �W         �W    �      �?N F�     �?N F�   �   ]  V  F ��-      j M Generic Library        � $                       �   %      �%         �%    �      �?N Z%     �?N Z%   �   ^  g  B ��;      k = Generic Library        � &                       �   %   �?N n�     �?N n�   �   a  ` ��)     l M Generic Library        �                        �         �         �    �   &   �?N ��     �?N ��   �   b  _  a ��;      m A Generic Library        �                        �         �1         �1    �   #   �?N N�     �?N N�   �     N  X ��-      n A Generic Library        � '                       �   (      �}         �}    �   $   �?N �1     �?N �1   �   l  h  [ ��-      o  Generic Library         & � +      �:         �:    �   p  	  L-U                          p M Generic Library       ! � )                       �   *      R�         R�    �   +   �?N ��     �?N ��   �   t    p ��;      q A Generic Library        � ,                       �   -      �b         �b    �   *   �?N �
     �?N �
   �   u  y  s ��-      r ] Generic Library        �                        �         r�         r�    �   ,   �?N Z     �?N Z   �   x  w  r ��M       s = Generic Library        �                        �   -   �?N 2�     �?N 2�   �   
  | ��)     t M Generic Library        � .                       �   /      ��         ��    �   )   �?N 2^     �?N 2^   �   }  ~  o ��;      u A Generic Library        � 0                       �         2[         2[    �   /   �?N v     �?N v   �   �  �  � ��-      v A Generic Library        �                        �         F-         F-    �   0   �?N ��     �?N ��   �   �  �  � ��-      w = Generic Library        �                        �   1   �?N F     �?N F   �   �  � ��)     x A Generic Library        �                        �   1      2^         2^    �   .   �?N r     �?N r   �   �   �  � ��-      y  Generic Library         & � 8      8         8    �   �  
  L-T                          z = Generic Library        �                        �   2   �?N �     �?N �   �   �  � ��)     { ] Generic Library        �                        �         �         �    �   3   �?N fq     �?N fq   �   �  �  � ��M       | A Generic Library        � 2                       �   3      RX         RX    �   4   �?N �\     �?N �\   �   �  �  � ��-      } A Generic Library        �                        �         "�         "�    �   5   �?N �~     �?N �~   �   �  �  � ��-      ~ A Generic Library        �                        �   5      ��         ��    �   6   �?N &�     �?N &�   �   �  �  � ��-       M Generic Library        � 4                       �   6      n�         n�    �   7   �?N v�     �?N v�   �   �  �  � ��;      � A Generic Library       ! �                        �   7      (         (    �   8   �?N �;     �?N �;   �   �   �  � ��-      �  Generic Library          � ;      ��         ��    �   �    L-S                          � A Generic Library        � 9                       �   :      �         �    �   ;   �?N ��     �?N ��   �   �  �  � ��-      � A Generic Library        �                        �         �         �    �   :   �?N 
�     �?N 
�   �     �  � ��-      � A Generic Library        �                        �         Z�         Z�    �   9   �?N jw     �?N jw   �   �  �  � ��-      � M Generic Library        � <                       �   =      �P         �P    �   >   �?N V�     �?N V�   �   �  �  � ��;      � G Generic Library       > � ?                       �   @      vD         vD    �   A      n         n    �   B      �T         �T    �   C      �H         �H    �   �  �  �  �  � ��3     �  Generic Library         ! � >      �         �    �   �    L-R                          � = Generic Library        �                        �   D   �?N ��     �?N ��   �   �  � ��)     � M Generic Library        �                        �         *�         *�    �   =   �?N ��     �?N ��   �     �  � ��;      � M Generic Library        � D                       �         b�         b�    �   <   �?N *,     �?N *,   �   �  �  � ��;      �  Generic Library         & � H      *�         *�    �   �    L-Q                          � = Generic Library        �                        �   E   �?N �S     �?N �S   �   �  � ��)     � M Generic Library       ! � F                       �   G      &@         &@    �   H   �?N ��     �?N ��   �   �  �  � ��;      � A Generic Library        �                        �   E      �y         �y    �   G   �?N Fk     �?N Fk   �      �  � ��-      � M Generic Library        � I                       �   J      ��         ��    �   F   �?N j�     �?N j�   �   �  �  � ��;      � A Generic Library        � K                       �         ��         ��    �   J   �?N 2�     �?N 2�   �   �  �  � ��-      � A Generic Library        �                        �         >�         >�    �   K   �?N ��     �?N ��   �   �  �  � ��-      � A Generic Library        � L                       �   M      �s         �s    �   I   �?N R�     �?N R�   �   �  �  � ��-      � = Generic Library        �                        �   M   �?N '     �?N '   �   �   � ��)     � ] Generic Library        �                        �         ^+         ^+    �   L   �?N �3     �?N �3   �   �  �  � ��M       � M Generic Library       & � N                       �   O      ��         ��    �   P   �?N �;     �?N �;   �   �  �  � ��;      � M Generic Library       ! � Q                       �   R                   �   O   �?N ��     �?N ��   �   �  �  � ��;      � M Generic Library       ! � S                       �   T      f\         f\    �   N   �?N 6k     �?N 6k   �   �  �  � ��;      �  Generic Library         + � P      �\         �\    �   �    L-P                          � = Generic Library        �                        �   U   �?N >�     �?N >�   �   �   � ��)     � = Generic Library        �                        �   V   �?N J�     �?N J�   �   �  � ��)     � A Generic Library        � W                       �         &�         &�    �   Q   �?N ��     �?N ��   �   �  �   � ��-      � A Generic Library        �                        �         ��         ��    �   W   �?N �     �?N �   �   �  �  � ��-      � A Generic Library        � V                       �   U      ��         ��    �   X   �?N �     �?N �   �   �  �  � ��-      � ] Generic Library        �                        �         �         �    �   Y   �?N �:     �?N �:   �        ��M       � A Generic Library        � X                       �         &�         &�    �   R   �?N ��     �?N ��   �   �  �  � ��-      � = Generic Library        �                        �   Z   �?N �7     �?N �7   �     	 ��)     � A Generic Library        � Y                       �   Z      V�         V�    �   T   �?N V�     �?N V�   �        ��-      � A Generic Library        � [                       �   \      V�         V�    �   S   �?N V�     �?N V�   �        � ��-      � = Generic Library        �                        �   \   �?N �7     �?N �7   �      ��)     � = Generic Library        � ]                       �   [   �?N "N     �?N "N   �       ��)     � ] Generic Library        �                        �         �         �    �   ]   �?N �:     �?N �:   �   !  �    ��M       �  Generic Library         + � `      �         �    �       L-O                          � M Generic Library       & � ^                       �   _      B         B    �   `   �?N �=     �?N �=   �   -     ��;      � M Generic Library       ! | a                       �   b      �w         �w    �   ^   �?N ��     �?N ��   �      "   ��;      �  Generic Library         ! r g      �         �    �   &    L-N                          � = Generic Library        u                        �   c   �?N (�     �?N (�   �   '  * ��)     � = Generic Library        s                        �   d   �?N �     �?N �   �   �   + ��)     � M Generic Library        q e                       �   f      Z�         Z�    �   g   �?N ��     �?N ��   �   /  4  & ��;      � M Generic Library        s d                       �   c      jF         jF    �   f   �?N Nl     �?N Nl   �   +  *  0 ��;      � = Generic Library        o                        �   h   �?N �f     �?N �f   �   1  2 ��)     � M Generic Library        o h                       �         >�         >�    �   e   �?N ��     �?N ��   �   2  )  , ��;      � = Generic Library        �                        �   i   �?N J�     �?N J�   �   �   8 ��)     � = Generic Library        �                        �   j   �?N �     �?N �   �   <  9 ��)     � A Generic Library        � j                       �   i      ��         ��    �   k   �?N �     �?N �   �   9  8  ; ��-      � A Generic Library        � k                       �         &�         &�    �   _   �?N ��     �?N ��   �   ;  ?   ��-      � A Generic Library         l                       �         &�         &�    �   b   �?N ��     �?N ��   �   E  �    ��-      � A Generic Library        ~                        �         ��         ��    �   l   �?N �     �?N �   �   F  B  E ��-      � M Generic Library       & a m                       �   n      ��         ��    �   o   �?N ��     �?N ��   �   c  Y  H ��;      � A Generic Library        y p                       �   q      Z_         Z_    �   a   �?N N�     �?N N�   �   I  K  J ��-      � = Generic Library        { r                       �   q   �?N ��     �?N ��   �   O  K ��)     � ] Generic Library        z                        �         ��         ��    �   r   �?N N�     �?N N�   �   �   P  O ��M       � = Generic Library        x                        �   p   �?N �      �?N �    �   R  U ��)     � = Generic Library        d                        �   s   �?N <&     �?N <&   �   �  Z ��)     � A Generic Library       ! e s                       �   t      ��         ��    �   n   �?N �$     �?N �$   �   X  [  \ ��-      � = Generic Library        ` u                       �   v   �?N vx     �?N vx   �   b  M ��)     � A Generic Library        ` v                       �         z�         z�    �   m   �?N �     �?N �   �   M  `  V ��-      � ] Generic Library        _                        �         ��         ��    �   u   �?N ڄ     �?N ڄ   �   f  �   b ��M       � ] Generic Library        f                        �         Z�         Z�    �   w   �?N >�     �?N >�   �   �  �   a ��M       � A Generic Library        W                        �   x      ��         ��    �   y   �?N ��     �?N ��   �   n  q  p ��-      � = Generic Library        Y                        �   x   �?N "9     �?N "9   �   v  q ��)     � M Generic Library        h w                       �   z      �4         �4    �   t   �?N ��     �?N ��   �   +  �  r ��;      � A Generic Library        [                        �         n�         n�    �   {   �?N �     �?N �   �   �   x  w ��-      � A Generic Library        Y y                       �   {      �V         �V    �   |   �?N �R     �?N �R   �   |  {  z ��-      �  Generic Library         ! Z |      �f         �f    �   z    L-L                          �  Generic Library         ! Q       b         b    �   ~    L-K                          � A Generic Library        P }                       �   ~      �V         �V    �      �?N �R     �?N �R   �   �  �  ~ ��-      � A Generic Library        R                        �   �      n�         n�    �   ~   �?N �     �?N �   �   �   �  � ��-      � = Generic Library        T                        �   �   �?N �     �?N �   �   �  � ��)     � = Generic Library        N                        �   �   �?N 6�     �?N 6�   �   �  � ��)     � A Generic Library        N �                       �         ��         ��    �   }   �?N ��     �?N ��   �   �  �  } ��-      �  Generic Library         ! H �      �@         �@    �   �    L-J                          � M Generic Library        G �                       �   �      �         �    �   �   �?N .�     �?N .�   �   �  �  � ��;      � = Generic Library        J �                       �   �   �?N ��     �?N ��   �   �  � ��)     � ] Generic Library        I                        �         ^          ^     �   �   �?N       �?N     �   �  �   � ��M       � M Generic Library        E �                       �   �      �'         �'    �   �   �?N B�     �?N B�   �   �  �  � ��;      � = Generic Library        G                        �   �   �?N 
0     �?N 
0   �   �  � ��)     � = Generic Library        E                        �   �   �?N f�     �?N f�   �   �  � ��)     �  Generic Library         + 7 �      t         t    �   �    L-I                          � M Generic Library       & 6 �                       �   �      �y         �y    �   �   �?N �}     �?N �}   �   �  �  � ��;      � M Generic Library       ! < �                       �   �      �l         �l    �   �   �?N q     �?N q   �   �  �  � ��;      � = Generic Library        A �                       �   �   �?N }     �?N }   �   �  � ��)     � A Generic Library        ?                        �   �      Z�         Z�    �   �   �?N 
�     �?N 
�   �   �  �  � ��-      � = Generic Library        <                        �   �   �?N �     �?N �   �   �  � ��)     � ] Generic Library        @                        �         �b         �b    �   �   �?N �^     �?N �^   �   �  �   � ��M       � A Generic Library        : �                       �   �      �|         �|    �   �   �?N �     �?N �   �   �  �  � ��-      � A Generic Library        9                        �         n�         n�    �   �   �?N �     �?N �   �   �  �   � ��-      � = Generic Library        7                        �   �   �?N       �?N     �   �   � ��)     � = Generic Library        5                        �   �   �?N 27     �?N 27   �   �  � ��)     � A Generic Library        5 �                       �   �      �         �    �   �   �?N &     �?N &   �   �  �  � ��-      � A Generic Library        4                        �   �      ��         ��    �   �   �?N ��     �?N ��   �   �  �  � ��-      � M Generic Library       ! 0                         �   �      �d         �d    �   �   �?N T�     �?N T�   �   ,  �  � ��;      �  Generic Library         + * �      ��         ��    �   �    L-H                          �  Generic Library         + ( �      ��         ��    �   �    L-G                          � M Generic Library        �                        �         �         �    �   (   �?N ��     �?N ��   �   �   j  h ��;      � = Generic Library        �                        �   '   �?N �     �?N �   �   i  f ��)     � M Generic Library        j                         �         �         �    �   �   �?N      �?N    �   �  ]  � ��;      �  Generic Library         + b o      �         �    �   H    L-M                          � M Generic Library       & ( �                       �   �      0h         0h    �   �   �?N <m     �?N <m   �   �  �  � ��;      � M Generic Library       ! % �                       �   �      *0         *0    �   �   �?N 65     �?N 65   �   �  �  � ��;      � = Generic Library        .                        �   �   �?N B9     �?N B9   �   �  � ��)     � A Generic Library        , �                       �   �      
[         
[    �   �   �?N >�     �?N >�   �   �  �  � ��-      � = Generic Library        , �                       �   �   �?N �u     �?N �u   �   �  � ��)     � ] Generic Library        +                        �         r�         r�    �   �   �?N ғ     �?N ғ   �   �  �   � ��M       � M Generic Library        '                        �         ��         ��    �   �   �?N n�     �?N n�   �   �  �  � ��;      � = Generic Library        k �                       �   z   �?N 
7     �?N 
7   �   �  � ��)     � = Generic Library        ( �                       �   �   �?N r     �?N r   �   �  �  ��)     � A Generic Library        " �                       �   �      �K         �K    �   �   �?N Ҵ     �?N Ҵ   �   �  �  � ��-      � = Generic Library        #                        �   �   �?N �     �?N �   �   �  � ��)     � M Generic Library        # �                       �                        �   �   �?N B�     �?N B�   �   �  �   � ��;      �  Generic Library         +  �      Ns         Ns    �   �    L-F                          � = Generic Library        !                        �   �   �?N ��     �?N ��   �   �   ��)     � M Generic Library       &  �                       �   �      N         N    �   �   �?N �M     �?N �M   �   �  �  � ��;      � M Generic Library       !  �                       �   �      &�         &�    �   �   �?N ֎     �?N ֎   �   �  �    ��;      � M Generic Library       !  �                       �   �      ��         ��    �   �   �?N ��     �?N ��   �     �  � ��;      � = Generic Library                                �   �      ��         ��    �      ��)     � = Generic Library                                �   �   �?N bq     �?N bq   �   �    ��)     � = Generic Library                                �   �   �?N �     �?N �   �      ��)     � A Generic Library         �                       �         
�         
�    �   �   �?N ��     �?N ��   �        ��-      � A Generic Library         �                       �   �      X�         X�    �   �   �?N ��     �?N ��   �        ��-      � A Generic Library                                �         �         �    �   �   �?N \�     �?N \�   �   	  �    ��-      � A Generic Library         �                       �         h�         h�    �   �   �?N HT     �?N HT   �     
   ��-       A Generic Library         �                       �   �      �-         �-    �   �   �?N ~�     �?N ~�   �       � ��-      = Generic Library                                �   �   �?N ��     �?N ��   �      ��)     M Generic Library                                �   �      �#         �#    �   �   �?N v�     �?N v�   �         ��;      = Generic Library                                �   �   �?N �     �?N �   �   "  # ��)     � �         �    �     !        �    �   �    �    �    �    �   �    �    �    �    �    �    �    �    �    z    r    �    l    e    ]    K    G   v    ~    �    �    �    �    �     !        �    �    �    �    �    �   �    �   �    �   �    �    �   �   �   �   r   l   h    e   \    X    Q    J    v   }    {    �   �    �    �    !     �    �   �   �    �   �   �    �    �   �    �    �   �    �   �   �    �    �    �    s    m    [    Y   P    N    �    x    �    �    �   �   �    #        �   �    �    �    �    �    �    �   �    �   �   �    �   �   �   �    �   �   w    �   m   g    ]   \   W    Q   L   I    u   }   {   �   �      F    P      F   O      F    E      G    H    	  G    M   
  H    J      H   I      K    L      L    M      M    O     N    O      P   Q      T    U      T   Y      T    R    S      U    ]      U   V      V    \      V   [      W    Z     X    Z      Y    Z      c    j      c   d      c    ^      d    i      d   f       e    f    !  f   g    "  h    i   #  i    m    $  j    n    %  j   k    &  k    l    '  n    �    (  n   �    )  p    t    *  p   q    +  p    o    ,  q    r    -  q   s    .  t    x    /  t   u    0  u    v    1  w    x   2  z    |    3  {    |   4  |        5  }    ~   6  ~       7      �   8  �    y    9  �    �    :  �   �    ;  �    �    <  �    �    =  �   �    >  �    �    ?  �    @  �   A  �   B  �   C  �    D  �    �    E  �    �   F  �    �    G  �   �    H  �    �    I  �    �    J  �   �    K  �    �    L  �    �    M  �   �    N  �    �    O  �   �    P  �    �    Q  �    �    R  �   �    S  �    �    T  �   �    U  �    �   V  �    �    W  �    �    X  �    �    Y  �    �    Z  �    �   [  �    �    \  �   �    ]  �    �    ^  �    �    _  �   �    `  �    �    a  �    �    b  �   �    c  �    �   d  �    �    e  �    �    f  �   �    g  �    �    h  �    �    i  �    �   j  �    �    k  �    �    l  �    �    m  �    �    n  �   �    o  �    �    p  �    �    q  �   �    r  �    �    s  �    �    t  �   �    u  �    �    v  �    �    w  �    �    x  �   �    y  �    �    z  �   �    {  �    �   |  �    �    }  �    �    ~  �   �      �    �    �  �   �    �  �    �    �  �    �    �  �   �    �  �    �    �  �    �    �  �    �    �  �   �    �  �    �    �  �   �    �  �    �    �  �    �    �  �   �    �  �    �    �  �    �   �  �    �   �  �    �    �  �    �   �  �    �    �  �    �   �  �    �   �  �    �    �  �    �    �  �   �    �  �    �    �    �  �    �    �  �   �    �  �    �   �  �    �    �  �    �    �  �    �    �  �    �    �  �   �    �  �    �    �  �    �    �  �   �    �  �    �    �  �    �    �  �   �    �  �        �  �   �    �  �    �   �  �    �    �  �    �    �  �    �    �         �        �       |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 7=� 1'� .1� �� ;.� �� �� .� :� 7� W.� 5��� ������ =�� =� � >�� ?@� C:� DW� AC� ;� E7� �� � Q>� � � ><� ?8� @E� A3� @2� 40� � � � D� Z?� PA� :� C-� :� �D� E&� \G� BH� YR� FI� ZJ� iZ� PK� eP� QL� dQ� eM� ce� iN� ni� �� q�� OT� :;� X]� g`� [^� c_� W� db� �d� fl� nj� m#� q� �  )� �i� "� �q� !� m� ��� 	5� y|� ru� �
� ��� zw� zc� {x� {�� 1^� s� ot� ~�� �n� �}� ��� ��� � � �� � ��� ��� �{� ��� ��� ��� ��� �� ������������������	��
���� ������������������������������������� ��!��"��#��$��%� &��'��(��)��*��+��,��-��.��/��0�� 1��2��3�4��5��6��7��8��9��:�;<��=��>m�?�@��A��B��C=mD@�E!F�G�H� IJKL	M
N@�OPQ
�RS�T.U=V=� W5X�YCZ@�[eG\WL]SN^3C_T3`u�a>
bN>cL.dm� eLRfT� gdThGPiG5jNFk.Bl3� m5?nU6ooSp6Iq><rC� s)dt�eu�Wv��w&oxS1y40z�){s�|,/}W)~d� e'�t��j"�J �����j�l�l�����z��,��������&�Z-��]�-��/�u��s��t��� �������������������������� �����f������ �����u�}���+�{w����� ��t�a���s��x�p|��n�&`�)� ����������[r����o�����������������������������Y\����������-X��� ����������������������� ����������� �������������������� �������������� ��������������������v�� ��������� ��� �	����
������� �!��$����*�Vc�,$�" ! ������%!%� () *	 ,	��
����$�%�$k#h#(00������������������	           ��������������������������������������������������������������)  	         �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �  �     �   �  �  x     �   � ! �  �       �  �  �     0  �    �    �  �           �    �     �  �  &  �    �  �  .  �    �  �  8  �     �  �  <  �    �  �  C  �    �  �  L  �    �  �  S  �     �  �  \  �     �  �  b  �    �  �  i  �    �  �  t  �     ~  �  {  �     f  �  �  �    l  �  �  �     r  �  �  �    H  � 0  E    F        � + 	 F    �   �  )  �     � � �  �  �    V  � !  M    �  	 � &  O   M        � !  G     �  	 �  �  �     d  �   G    H        �   G    �   �   H   I        �   H    J       
 �   I     �     �  �     %    J     �    �  �     3    L     �     L    �     K    L        !  M     �    �  �       +  F     �   	 	 N     �   
 �  s     �   �� �  m     �            �     �  [     �   +  O     �     K     �   &  O     �     Q    �     Q     �     P     �     P   Q        ��  P     �     Y    �   & �  T     �   & �  R     �    �  ]     �    �  V     �   & �  S       ��! �  T     �    ! �  T    �   ! �  U    �   "! �  U     �   # �  U     �   $ �  V    \        ��&  W     �   '  W    Z       ( �  X    Z        )!  Y     �   ��+   Y    Z        ,! 1  �     �   - �  X     �   .    � � �   ��0 �  [     �   1 	   � � �   2 �  \    �   3 �  \     �   4 �  V    �   5& 	   � �   ��7    � � �   8 �  ]    �   9& �  ^    c        :    � � �   ;    � � �   < �  ]     �   =    � � �   > �    � � �   ? �    � � �   @ �    � � �   A �    � � �   B! �  j     �   C �    � � �   D �    � � �   E    � � �   F �  i     �   G! �  d     �   H! �  c     �   I �  d     �   J �  g     �   K �  e    �   L �  e     �   M �  h     �   N �  m    �   O �  e     �    P �    � � �   Q �    � � �   R �  f     �   S �  f   g       ! T �  f     �    ��V �  h    i      " W    � � �   X �  m     �  # Y �  d    �   Z �    � � �   [ �  n     �  $ \! �  c    �   ] �  i     �  # ^ �  j     �  $ _ �  l    �   ` �  k     �  % a �  k    l       & b �  l     �   c �    � � �   d �    � � �   e �    � � �   f �  �     �  ' g �  j    �  % h �  �    n      ( i �    � � �   j �  �    �   ��l �  n     �  ' m �    � �   n �    � � �   o! �  t     �  ) p& �  p    o       + q �    � � �   r �  r     �  , s �  q     �  * t! �  p     �  ) u �  q     �  , ��w �  r    �   x �  r     �   y �  q    �  - z �    � ��   { �    � � �   | �  s     �  - } �  t     �  . ~ �  t    �  / ! �  p    �  * � �    � � �   ��� �  u    �   � �  v    �   � �  u     �  / � �    � � �   � �  v    u       0 � �  v       � �    � ��   � �    � �   ��� �  x   w       1 � �    � � �   � �  x     �  . � �  }    ~      5 � �  z    |       2 � �  z       � �  {    |      3 � �  w     �   � �  {      �& �  �    y       8 �    � � �   � k  �     �   � �        4 � �  {     
  ��� �  }      � �  }     ,  �    � � �   � �    � 
  � �       6 � �  ~      6 � �  ~       �! �  �     7 �! �        7 � �    � � ,  � �  |      4 ��� �    � � �   � �     �   � �  �      9 � �  �    �       ; � �    �   � �  �      9 � �  �      ��� �  �      � �  �       � �  �      : � �    	   � �    �   � �  �     : ���! �  �    �       > � �      � �  �     = �C �  �       C �> �  �      B �> �  �      A �> �  �      @ � �  �      < � �  �      < � �  �    5  ��� �  �    1  � �  �    �       D � �      �> �  �       ? � �      � �      � �  �      = � �    	  �! �  �     " F �& �  �    �       H � �  �     *  �! �  �     " F � �  �    �      E � �  �     #  � �    %&  � �  �     ! G ��� �  �     ( I �! �  �    ! G � �    #$  � �  �     ( I � �  �    )  � �  �    +  � �  �     ' J � �    )$S  � �  �    �       K � �  �     -  � �    +A  � �  �    ' J � �    -.   � �  �    �       L ��� �  �     / M � �    &>0  � �  �    2  �& �  �     7 N �+ �  �    �       P � �  �     4  �! �  �    9 R �& �  �     6 O �! �  �     8 Q �! �  �    : T �! �  �     < S �& �  �    6 O �& �  �     7 N �! �  �     < S � �  �    / M � �    2A@  � �    4.N  ��� �  �    �      U � �  �    �       V � �    *   � �  �    �       X � �  �     Z  � �    1  �! �  �     9 R � �  �     8 Q � �  �    X  ��� �    3  � �    5  ��� �    GF \   �  �    �       [  �  �    �       ] �� �  �    �       Y  �    JG \  �  �     P   �    ETK   �  �    O   �    IW�  	 �  �     L Z 
 �    MaQ   �  �     ; T  �  �    L Z  �  �    J \  �    ;: T �� �  �     M  �� �    PK?  �� �    HUY   �    O�R   �  �     F \  �  �     I   �    XSR  ! �  �     � _ & ~  �     � ^ + �  �    �       `            �  �     � b  �     & �  �    � _  ! }  �     � a ! �  �     E  "!   �    � b # �     $ �     % �     &! s  �    �       g ' v  �       ��) r  �    }  * v  �    �      c + t  �    �       d , q  �     | e -& �  �     � ^ . �    kcT  / r  �     | e 0 u  �     y f 1 p  �     x  2 p  �    �       h 3 �    l^_  4 t  �    y f 5 �    miW  6 y    pn p ��8 �  �    �      i 9 �  �    �       j :+    � �   ; �  �    �       k < �  �     q  = �    VCU  > �    qba  ? �  �    m  @ �    ZND  ��B �  �    k  C �    rY^  ��E �  �    �       l F   �     j  G }    h[i  H+ c  �    �       o I z  �     p p J! {  �     � a K |  �   �       q L y    e\c  M a  �    �       v N     j]b  O |  �    �       r P }  �    h  ��R y  �     e  S p    xo]  T {    f_g  U y  �     n p V! b  �     � m W r    }u\  X! f  �     � s Y& d  �    � n Z e  �     � s [! h  �    � t \& g  �     � n ] m  �    �  ^ 	 N     �   ��` c  �    �  a h  �     � w b a  �    �       u c& b  �     � m d t    ~gs  e v    t[  f `  �     �  ��h :     i �  �     �   j     �� b k =     l! �    �� _ m �    d>C  n X  �     �  o e    wo�  p Y  �     � y q Z  �    �      x r! j  �     � t s H    ��{  t J    ���  u F    ��`  v Z  �     �  w ]  �     � { x ^  �    �  ��z! [  �    �       | { \  �    � { | Z  �     � y } P  �     � } ~! R  �    �         L    ���  � Q  �     � } � <     � U  �     �  ��� Q  �    �  � T  �     � ~ � U  �   �       � � O    �`�  � 9     � O  �     �  � O  �    �       � � S    ���  � S  �    � ~ � \    ���  � G  �     � � �! I  �    �       � � Q    ���  � K  �     � � � K  �    �       � ��� J  �     �  � H  �     � � � Z    ���  � U    �{�  � J  �    � � � H  �   �       � � F  �    �       � � H  �     �  � ^    ���  � F  �     �  �& 2  �      � �& 9  �     � �+ 8  �    �       � � X    ���  �! =  �     
 � ��� �  �    =  �& 7  �      � � B  �    �      � � g  �       � B  �    �       � � �  �    �       W �! A  �     � � � A  �     �  � �    ?@=  � =  �    � � � =  �     � � � �    � � �   � �    QDB  � :  �     �  � @  �       � m    �t�  �! <  �     
 � � =  �     �  � ;  �    �       � � e  �     �  � g    vu  � l  �    �       � � 5  �     �  � 6  �     �  � 7  �   �       � � 8  �    �      � � �    � � �   � 6  �    �       � � )  �    �       � �     ��    �! 6  �     � � �! 3  �    � � �! +    �� � � (    �� � � 1    ��	   �+ )  �     � � � /    ���  � $    ���  � .    ���  � &    ���  � ,    ���  � (    ���  � k    	��   � *    ���  � "    ���  � "    �� � �! .  �     � � �& )  �     � � �+ +  �     � � �& +  �    � � � �  �     B  �! &  �     � � �& '  �     � � �! (  �    � � �+ *  �     �� � � /  �    �      � � 8    ���  � /  �     �  � -  �    �       � � -  �    �       � � b    �z�  � *  �    �  � ,  �     �  � 6    ���  � 5    ���  � `    ��v  � =    ���  � @    ��  �! ?  �    � � � (  �     �  � l  �     � z � :    ���  � k  �    � z � #  �     � � �! $  �     � � � %  �   �       � � <    ���  � h    �� w � $  �    �       � �+   �    �       � � A    ���  � C    ���  �& >  �      � � $  �     �  �&   �     � � �&   �    � � �!   �     � � �!   �    � � � "  �     �  �&   �     � � �!   �    � � �!        � �  &   �     � � !     �� � !   �     � �    �     �     �    �      �    �    �       �      ���      �    �      � �   	   �     �  
   �    �     �    �       � !   �     � �       ���     �    �       �      ���   "  �     � �     �        ���     �     � �      ��       ���     �     � �      ���          � !     �� �          �    �     �                      �      ���          �            !      �  "       �  #        � $     ��  %       & c    ��w  '    �   (       ) i    sz�  * 	    �  + i  �     � w ,     �  -! e    �� s .    �   /    �              A      B     C     D     E   E  L-Z E  R  L-Y R  S  L-X S  ^  L-V ^ 	 o  L-U o 
 y  L-T y  �  L-S �  �  L-R �  �  L-Q �  �  L-P �  �  L-O �  �  L-N �  �  L-M �  �  L-L �  �  L-K �  �  L-J �  �  L-I �  �  L-H �  �  L-G �  �  L-F � ��                               	   
                            
   	                + V�     �An                                                         