      Generic Library                                   �        Set                           Generic Library                                  �    	     Reset                       �� < Generic Library                                �          �         �    �      �?N �     �?N �   �           ��(      < Generic Library                                �         �         �    �      �?N �     �?N �   �   	        ��(       Generic Library         2        H�         H�    �        Q                              Generic Library         2        ��         ��    �   
     No Q                                                                                   
                      	   
  	                 	          
         '           '                                ' 	         2            "           	         
   
 2            "                        '            	                 	              	             
   ������          Reset  ��    Set      Q     No Q                  2 _ ��     �?N                                                          