      Generic Library                                   �         .�         .�    �         ޢ         ޢ    �         ��         ��    �         A                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       B                             Generic Library          	                        �   	      .�         .�    �   
      ޢ         ޢ    �         ��         ��    �       C                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       D                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       E                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       F                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       G                             Generic Library                                  �         .�         .�    �         ޢ         ޢ    �         ��         ��    �       H                             Generic Library                                   �   !      .�         .�    �   "      ޢ         ޢ    �   #      ��         ��    �       I                           	  Generic Library           $                       �   %      .�         .�    �   &      ޢ         ޢ    �   '      ��         ��    �   	  	  J                           
  Generic Library          " (                       �   )      .�         .�    �   *      ޢ         ޢ    �   +      ��         ��    �   
  
  K                             Generic Library          % ,                       �   -      .�         .�    �   .      ޢ         ޢ    �   /      ��         ��    �       L                             Generic Library          ( 0                       �   1      .�         .�    �   2      ޢ         ޢ    �   3      ��         ��    �       M                             Generic Library          + 4                       �   5      .�         .�    �   6      ޢ         ޢ    �   7      ��         ��    �       N                             Generic Library          . 8                       �   9      .�         .�    �   :      ޢ         ޢ    �   ;      ��         ��    �   '    O                             Generic Library          1 <                       �   =      .�         .�    �   >      ޢ         ޢ    �   ?      ��         ��    �       P                             Generic Library          4 @                       �   A      .�         .�    �   B      ޢ         ޢ    �   C      ��         ��    �       Ctrl                          Generic Library#  	              v�         v�    �         �G         �G    �         *G         *G    �         �F         �F    �         �         �    �         �         �    �         ��         ��    �         �         �    �         h         h    �   	      ��         ��    �   
      n�         n�    �         ��         ��    �         �         �    �         d�         d�    �         8�         8�    �         JE         JE    �         �D         �D    �         ��         ��    �         ��         ��    �         �         �    �         
�         
�    �         �x         �x    �         D�         D�    �         �S         �S    �         �         �    �         Pf         Pf    �         J�         J�    �         S         S    �         4�         4�    �         @r         @r    �         ƫ         ƫ    �          �          �    �   @      �         �    �   A      |�         |�    �   B      �         �    �   D      f�         f�    �   E      2�         2�    �   F      Pq         Pq    �   G      ��         ��    �                           7   )  ��  v��O
 MUX3X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX3X4.CKT
 MUX3X4.CKTA � �o    B � �o   C � �o   D � �o   E � �o   F � �o   G � �o   H � �o  	 Ctrl  �o   
 Out0  �o    ������������������������������������������������������������������������������ �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  ��! ��" ��# ��$ ��% ��  �� ��* ��+ ��, ��- ��. ��     Generic Library       G         �6         �6    �         н         н    �         ��         ��    �         ��         ��    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �   	      8�         8�    �   
                   �         �         �    �         ��         ��    �         �         �    �         ��         ��    �         ��         ��    �         l�         l�    �         ��         ��    �         ��         ��    �         H�         H�    �         ��         ��    �         �         �    �                    ��  6��O
 MUX2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX2X4.CKT
 MUX2X4.CKTCtrl  W�    A rl  W�   B rl  W�   C rl  W�
   D rl  W�   Z rl  W�    �������������������������������������������� �� ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
     Generic Library	                vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �   	      .I         .I    �   
      ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	               vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	       % 
 	      vw         vw    �   
      %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library               ,          ,    �         <*         <*    �         �)         �)    �         �)         �)    �          ��                          ������������          ��        ��        ��        ��        ��        ��        ��        �� 	          ��   	           
                                 �� 
      ��       ��       ��       ��       ��       ��       ��                                        ��        ��        ��       ��       ��    Generic Library       G !        �6         �6    �         н         н    �         ��         ��    �         ��         ��    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �         8�         8�    �                      �         �         �    �          ��         ��    �   !      �         �    �   "      ��         ��    �   #      ��         ��    �   $      l�         l�    �   %      ��         ��    �   &      ��         ��    �   '      H�         H�    �   (      ��         ��    �   )      �         �    �                    ��  6��O
 MUX2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX2X4.CKT
 MUX2X4.CKTCtrl  W�    A rl  W�   B rl  W�   C rl  W�
   D rl  W�   Z rl  W�    �������������������������������������������� �� ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
     Generic Library	                vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �   	      .I         .I    �   
      ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	               vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	       % 
 	      vw         vw    �   
      %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library               ,          ,    �         <*         <*    �         �)         �)    �         �)         �)    �          ��                          ������������          ��        ��        ��        ��        ��        ��        ��        �� 	          ��   	           
                                 �� 
      ��       ��       ��       ��       ��       ��       ��                                        ��        ��        ��       ��       ��    Generic Library	       P        &         &    �         �         �    �         ʵ         ʵ    �         �         �    �   &                     �   '      �         �    �   (      �         �    �   )      �          �     �   *      �         �    �   +      �         �    �   ,      d�         d�    �   -      �0         �0    �   .      6         6    �               ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_�;_    A1 ;_�;_   B0 ;_�;_   B1 ;_�;_   Ctrl0 �;_   Z0 l0 �;_    Z1 l0 �;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��  �������������������� ` Generic Library      ? '        ZU         ZU    �         ��         ��    �   *      �k         �k    �          Ϊ         Ϊ    �         T�         T�    �   *      ��         ��    �   +  ,  .     ��	                                    ` Generic Library       B '        �         �    �         ��         ��    �          p         p    �         ̃         ̃    �   +   ,     ��                          / /         ��             �� !          ��         ��        ��        ��        ��        ��        ��  	     	 ��  
     
 ��        �� 	       �� 
       ��        ��        ��        ��        ��                                             ��       ��       ��       ��       ��       ��       ��      	 ��      
 ��       ��        ��  !     ��  "     ��  #     ��  $     ��  %     ��  &         '        (        )        *     �� " +      ��   ,     ��  -     ��  .     ��    Generic Library#  	      )        v�         v�    �   !      �G         �G    �   "      *G         *G    �   #      �F         �F    �   $      �         �    �   %      �         �    �   &      ��         ��    �   '      �         �    �   (      h         h    �   )      ��         ��    �   *      n�         n�    �   +      ��         ��    �   ,      �         �    �   -      d�         d�    �   .      8�         8�    �   /      JE         JE    �   0      �D         �D    �   1      ��         ��    �   2      ��         ��    �   3      �         �    �   4      
�         
�    �   5      �x         �x    �   6      D�         D�    �   7      �S         �S    �   8      �         �    �   9      Pf         Pf    �   :      J�         J�    �   ;      S         S    �   <      4�         4�    �   =      @r         @r    �   >      ƫ         ƫ    �   ?       �          �    �   @      �         �    �   A      |�         |�    �   B      �         �    �   H      f�         f�    �   I      2�         2�    �   J      Pq         Pq    �   K      ��         ��    �                  !   8   #   5   +  ��  v��O
 MUX3X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX3X4.CKT
 MUX3X4.CKTA t0  �o    B t0  �o   C t0  �o   D t0  �o   E t0  �o   F t0  �o   G t0  �o   H t0  �o  	 Ctrl  �o   
 Out0  �o    ������������������������������������������������������������������������������ �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  ��! ��" ��# ��$ ��% ��  �� ��* ��+ ��, ��- ��. ��     Generic Library       G         �6         �6    �         н         н    �         ��         ��    �         ��         ��    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �   	      8�         8�    �   
                   �         �         �    �         ��         ��    �         �         �    �         ��         ��    �         ��         ��    �         l�         l�    �         ��         ��    �         ��         ��    �         H�         H�    �         ��         ��    �         �         �    �                    ��  6��O
 MUX2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX2X4.CKT
 MUX2X4.CKTCtrl  W�    A rl  W�   B rl  W�   C rl  W�
   D rl  W�   Z rl  W�    �������������������������������������������� �� ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
     Generic Library	                vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �   	      .I         .I    �   
      ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	               vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	       % 
 	      vw         vw    �   
      %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library               ,          ,    �         <*         <*    �         �)         �)    �         �)         �)    �          ��                          ������������          ��        ��        ��        ��        ��        ��        ��        �� 	          ��   	           
                                 �� 
      ��       ��       ��       ��       ��       ��       ��                                        ��        ��        ��       ��       ��    Generic Library       G !        �6         �6    �         н         н    �         ��         ��    �         ��         ��    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �         8�         8�    �                      �         �         �    �          ��         ��    �   !      �         �    �   "      ��         ��    �   #      ��         ��    �   $      l�         l�    �   %      ��         ��    �   &      ��         ��    �   '      H�         H�    �   (      ��         ��    �   )      �         �    �                    ��  6��O
 MUX2X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX2X4.CKT
 MUX2X4.CKTCtrl  W�    A rl  W�   B rl  W�   C rl  W�
   D rl  W�   Z rl  W�    �������������������������������������������� �� ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
     Generic Library	                vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �   	      .I         .I    �   
      ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	               vw         vw    �         %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��    Generic Library	       % 
 	      vw         vw    �   
      %         %    �         ��         ��    �         ��         ��    �         �f         �f    �         �         �    �         �         �    �         J�         J�    �         ̃         ̃    �         .I         .I    �         ��         ��    �         H�         H�    �         8�         8�    �              ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_;_    A1 ;_;_   B0 ;_;_   B1 ;_;_   Ctrl0 ;_   Z0 l0 ;_    Z1 l0 ;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library               ,          ,    �         <*         <*    �         �)         �)    �         �)         �)    �          ��                          ������������          ��        ��        ��        ��        ��        ��        ��        �� 	          ��   	           
                                 �� 
      ��       ��       ��       ��       ��       ��       ��                                        ��        ��        ��       ��       ��    Generic Library	       P        &         &    �         �         �    �         ʵ         ʵ    �         �         �    �   &                     �   '      �         �    �   (      �         �    �   )      �          �     �   *      �         �    �   +      �         �    �   ,      d�         d�    �   -      �0         �0    �   .      6         6    �               ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 ;_�;_    A1 ;_�;_   B0 ;_�;_   B1 ;_�;_   Ctrl0 �;_   Z0 l0 �;_    Z1 l0 �;_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��  �������������������� ` Generic Library      ? '        ZU         ZU    �         ��         ��    �   *      �k         �k    �          Ϊ         Ϊ    �         T�         T�    �   *      ��         ��    �   +  ,  .     ��	                                    ` Generic Library       B '        �         �    �         ��         ��    �          p         p    �         ̃         ̃    �   +   ,     ��                          / /         ��             �� !          ��         ��        ��        ��        ��        ��        ��  	     	 ��  
     
 ��        �� 	       �� 
       ��        ��        ��        ��        ��                                             ��       ��       ��       ��       ��       ��       ��      	 ��      
 ��       ��        ��  !     ��  "     ��  #     ��  $     ��  %     ��  &         '        (        )        *     �� " +      ��   ,     ��  -     ��  .     ��    Generic Library	       +  D      n�         n�    �   E      $�         $�    �   F      ��         ��    �   G      ��         ��    �   H      J         J    �   I      h         h    �   J      �         �    �   K      D�         D�    �   C                   �   L      ��         ��    �   M      ��         ��    �   N                     �   O      `         `    �   *   %      (  ��  膙O
 MUX1X4.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X4.CKT
 MUX1X4.CKTA t0  �o    B t0  �o   Ctrl  �o   Z rl  �o    ��������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� ��  ����  Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 s W�    A1 s W�   B0 s W�   B1 s W�   Ctrl0 W�   Z0 l0 W�    Z1 l0 W�   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 <_<_    A1 <_<_   B0 <_<_   B1 <_<_   Ctrl0 <_   Z0 l0 <_    Z1 l0 <_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          �� ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                 ��     ��         ��       ��        ��       ��       ��       ��       ��          ��     	      ��   
     ��        ��       ��   ` Generic Library       5 @      �         �    �   A      �/         �/    �   B      �4         �4    �   C      ֥         ֥    �   @      ��         ��    �   A      ��         ��    �   B      ��         ��    �   C      J�         J�    �   4  3  2  "     ��
                                             ` Generic Library        5 @      r�         r�    �   A      ��         ��    �   B      �         �    �   @      Z9         Z9    �   A      8/         8/    �   B      ��         ��    �   $   ,   -   6  ��                                     Generic Library         3  L                       �   M      	         	    �   N      �         �    �   O      ڻ         ڻ    �   (     Z                            P P                                                                                  	       	 
       
                                                                                                                                                                                         !        "        #        $  	       %  	      &  	      '  	      (  
       )  
     	 *  
     
 +  
      ,         -        .        /        0         1        2        3        4         5        6        7        8         9        :        ;        <         =        >        ?        @              A       !   ! B       "   " C        D          E        F        G        H         I        J        K        L          M        N        O        ; ;   )    *  & %  & +   #  / 5  1 7  1 /  2 - 	 3 , 
 4 $  0 /  6 0  " .   .  '    8    !  9     9   :  : ;  ;   <   = <   =  
 >  > ?  ?   @   A @  	 A    B ! B C " C  # D  $ E D %   E & F  ' G F (  G ) H  * I H +  I , J  - J K .  K / L  0 L M 1  M 2  N 3 O N 4 O  5 P  6 P Q 7  Q 8  R 9 S R : S  U T            %                (        
       +   	 
           .               1               2               7               8                    ! " # 	     	       $ % & ' 
  #  
       ( ) * +   &         , - . /   )         0 1 2 3   ,         4 5 6 7   1       8 9 : ;   2         < = > ?   5             @ A B C   	       #         
      &              )   	 
          ,              /              4              5              :       +         C  "         D E F G   +       "    ! " #   ,        $ % & '   -        ( ) * +   .        , - . /   /        0 1 2 3    0       4 5 6 7 !  0        4 5 6 7 "  8        C #  2        < = > ? $  5       
  @ % +         H I J K & "        H I J K '  /         8 9 : ; ( 3              L M N O ) " 	          D E F G * +          D E F G + " +         H I J K ,  6      	  A -  7        B . + 8       C /  3        @ A B 0  5       @ A B 1         @ A B 2  7        B 3  6      	  A 4  5       
  @ 5  3        @ A B 6  5         @ A B 7          @ A B 8  1        8 9 : ; 9  ,       4 5 6 7 :  )       0 1 2 3 ;  /       0 1 2 3 <  .       , - . / =  &       , - . / >  #       ( ) * + ?  -       ( ) * + @  ,       $ % & ' A          $ % & ' B        !    ! " # C  +    ! "    ! " # D  	    # $       E      $ %       F  
    & '      G      ' (      H      ) *   	 
  I  
    * +   	 
  J      , -      K      - .      L      / 0      M      0 1      N      2 3      O      3 4      P      5 6      Q      6 7      R      8 9      S      9 :      ��   ��       A      B     C     D     E     F     G     H     I  	 	  J 	 
 
  K 
    L     M     N     O     P     Ctrl     Z                                 	 	  
 
                         ( ��      �An                                                         