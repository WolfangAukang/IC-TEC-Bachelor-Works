      Generic Library                                   �         A                             Generic Library          
                        �        B                             Generic Library                                  �        Ctrl                          Generic Library         %                         �        Z                             = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;                                                                                                               	    
  	                   	            	              %                 
                                         	         	         
   �� $                        	                                                                                                         A      B     Ctrl     Z  ��                 L ��       �An                                                         