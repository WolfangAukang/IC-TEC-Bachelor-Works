      Generic Library         6  	      �         �    �          C                              Generic Library         6  
      3         3    �        U                              Generic Library         6        >�         >�    �        D                              Generic Library         6 "       ��         ��    �        T                              Generic Library                                   �        A0                            Generic Library                                  �        A1                           = Generic Library       
                        �      �?N �l     �?N �l   �       ��)      = Generic Library       
                         �      �?N �l     �?N �l   �     	  ��)      A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �   
        ��-      	 A Generic Library       %                          �         �#         �#    �      �?N �#     �?N �#   �           ��-      
 A Generic Library       %                         �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       %                           �         �#         �#    �      �?N �#     �?N �#   �           ��-       A Generic Library       /                         �         �#         �#    �   	   �?N �#     �?N �#   �   '   (     ��-       A Generic Library       /                         �         �#         �#    �   
   �?N �#     �?N �#   �         !  ��-       A Generic Library       /                         �         �#         �#    �      �?N �#     �?N �#   �   %        ��-       A Generic Library       / !                        �         �#         �#    �      �?N �#     �?N �#   �   #   $     ��-        Generic Library          $                        �   "     Hab                                  	                     
                 	             
               	          
                                    	           
                              ' '             !               $  " & 	 &   
           '   (   %   #   /  ) 
  	 )     +    +  0 *  *   -   . 2  ,      . /  /   , 0   0  ! 1  " + 1 # - 2 $ 2  % 3  & ) 3 5 4   6           	  6          
  6            6 #                                                  
            
           	            
 %            %           *            %   	           %   	    !    *   	         %   
     $    %   
    %    * "           % !            % #          *   
         /            ,      
    4 #            /           ,       
    4            /           ,           4          	               , $    	     ! 4          
 "  %          # / "          $ / $         % /           & , %     	   ' /           ( /          )        &   * # !         +        "   , #          - " #     #   . "         /           0 #            1      ! "   2 "     #  $   3      % &   ��           C      U     D     T     A0     A1     Hab                            L ��       �An                                                         