      Generic Library                                   �         ܳ         ܳ    �         ��         ��    �         <�         <�    �         A                             Generic Library                                  �         ��         ��    �         D�         D�    �         ��         ��    �       B                             Generic Library                �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �   	      X|         X|    �   
      �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0  a�G    A1  a�G   B0  a�G   B1  a�G   Ctrl0 a�G   Z0 l0 a�G    Z1 l0 a�G   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library               ��         ��    �         2          2     �          �         �    �         ��         ��    �   
  	     ��                           ` Generic Library              �         �    �         2�         2�    �         ��         ��    �         ��         ��    �          ��                           ` Generic Library               ��         ��    �         ��         ��    �         ��         ��    �         Z�         Z�    �          
�         
�    �         ��         ��    �         j�         j�    �         �         �    �   !        ��                                  ` Generic Library       	       f�         f�    �         ��         ��    �         2�         2�    �         ��         ��    �         ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �           ��                                   Generic Library               �          �     �                        �         8�         8�    �         ��         ��    �         �         �    �         X|         X|    �         �w         �w    �                      ��  ���O
 MUX1X2.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X2.CKT
 MUX1X2.CKTA0 <_z<_    A1 <_z<_   B0 <_z<_   B1 <_z<_   Ctrl0 z<_   Z0 l0 z<_    Z1 l0 z<_   ��������������  �� �� �� �� �� �� ��
  ��������������  Generic Library                ��         ��    �         
         
    �         �         �    �         8�         8�    �         	     ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA �s W�    B �s W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��     Generic Library               ��         ��    �         
         
    �         �         �    �         8�         8�    �              ��  6�O
 MUX1X1.CKT2 C:\USERS\KIRSTEIN\AKW\ISEMES~1\B2LOGIC3\MUX1X1.CKT
 MUX1X1.CKTA rl  W�    B rl  W�   Ctrl  W�   Z rl  W�    ��������  �� �� �� ��  �������� = Generic Library                               �      �?N 8v     �?N 8v   �     	  ��)      A Generic Library                                 �         �Q         �Q    �      �?N >Q     �?N >Q   �           ��-       A Generic Library        
                        �         �Q         �Q    �      �?N >Q     �?N >Q   �            ��-       M Generic Library                                �         JG         JG    �      �?N �F     �?N �F   �           ��;           ��         ��        ��                                           ��   ��     ��         ��        ��       ��       ��              ��         ��   ` Generic Library              ��         ��    �         
�         
�    �         ��         ��    �         j�         j�    �          ��                          	 ` Generic Library              �         �    �         6�         6�    �         ��         ��    �         ��         ��    �          ��                          
  Generic Library                                  �        Ctrl                         ` Generic Library       $  	      F�         F�    �   
      b�         b�    �   	      �         �    �   
      ��         ��    �         #  ��                           ` Generic Library       $        ��         ��    �         ��         ��    �         ��         ��    �         V�         V�    �         %  ��                           ` Generic Library       '  	      :�         :�    �   
      V�         V�    �         �         �    �         ��         ��    �   	      f�         f�    �   
      �         �    �         ��         ��    �         v�         v�    �   "   %   &  ��                                   Generic Library         *  	                       �   
      �         �    �         ��         ��    �         N�         N�    �   &     Z                                                                                                            
       	          
                             	   
         !               	   
                " # ( &                         	                                                                           
         $              	  $            
 	            
                                                    	     
                       	 
                                  	               	                   $                $                                      
      	                                                                 	           !              " '          	 
 # '          	 
 ��% '               & *              	 
   ��           A      B   
  Ctrl 
    Z                   E �y       �An                                                         